
// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype.sv"
`define PATNUM 100000
`define SEED 45
`define CYCLE 15


program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
#];GNMQN206Kf,4F;4_bK6QSZ\^1RG0F,E\B.177^PMWSQ7@A8927)H](YTTQRa=
eS9RS<cJ=_b07dZW_S6.=[F3DC6<a).ILU_3Y?cBRWR9TEg\H2[P_e6_J4BOZ_A1
7+VVS9L]<bYNSTF,[O2R[9?8NCDTZT5P6PQQR@:cWZ1EQCOCDALf@E<&4UM05gT#
&0A1H/f8UAMSeW;eY8X[fEP)=A](f;M)@T5#:7P]QL499@9.=825^:?]TKLMWV1<
<PLX:eGD(_8UB^TS5WQ)a:#d]gWF7VB6(APEI?3IKV-\_Ee5-R#9S=@(OIK,TN\_
3#ZAG:\]OS<?3B[,5?X6YX3^)XeCAR96f>X<USFdB&T8Ke<6+W)0Xe4FP1O<fOEP
5aW_;(aG6,5/?SU/VN+A43LUZS7XO7?7DTSa_;bQd]4PWFN7c,;CT-A[a:N0F7.0
((I[QZQGKWa6>MC691B4dV.UD]B,D;dOJ&Q=gK3CQ,6;0WfX?2PU_;N_1,Y&W5]1
G7GMdfO+I/GJN@^Q>E:M?N]U(2?\9\((SLb:G#?,D83>_WUPPK/[54#eKN]FQe/-
8d6G7,^#-DWO+9()M8c54/SeXDHf.bU752IPKfR;/CN^?/,@01X-3#;N/-TS?MR^
5@\;CdY1cY3a\(.=MLJ/BN0g.:)f#[/3g)f9B?+/_c?gSWO)_]VN>@AXR^7,,)&d
.>5:cA(,F-J:g,Q5-5CSba@,T#CF]d]0_:2H;SA)3G^Yd>g0^0<:D8^F.]U1-Jac
H^#)?>C[\9T&PRc>6PZ8,^#9U7[a@e]E=\W>30,4-V?[gSeU^?MIcX^+GdUMS/WZ
?=@BHIN1S6-3B;RJ(2@E=S:COJ41?c?K_La6fQ4D4Y-dS2Xb5g^4[RWaZ4da1\I?
KW14eYIGD8?[^;>ZSE\+BaS^DDS(R[&?b4Z#PWe;B3gg#\+GH18S6]M_6G\=T:DJ
+K8F69CE@Ve=6BF<HcQ@V;B\::4^dVBHBWGET[+[&\=,&63<]U)EW?Y&65W9P4eM
8_:g/@O2G[9bg;(^3V>S>#d3bXHS]7e.XAIDW#M4V:/UVSSC59BJ]5aEY=GF>Hba
]DHW.1-8>.A]d;=[;S&ODCOE?\eJ7;AC>\JJ,ag\VTYDX-D.3f47@GN861]f,Gg6
O05;A_Pa@56EHBEF<Y]GFY/5PLOXCdU2VD-PI<WYDK[bP1MB@/a@X&W/U,>FSV,E
L.>+:Wg[8GDVTLC^I9(-E&Ef_3ULbVI/((>SGLBdUFJ0#)4A@R3.8@[R211cdTMI
ND6>bS\e-c6[R\#H^VZ,acENG4M84aTURA<QObF.46GD4FIE#c8AO>MbOM8&-V[,
DX\5\^Y-cEVf4/)S\K]XdMfH=2<NcZGSUOa:P+W?EWFKR+GDX7f5dA7Vc?]9b=[A
.N5\@^=_1F6;67fC&8VW:J4J9V5FV+Mg\@8F[2J=H4F&f1D?bVLd:P?TcQZ;,GFX
92QV^?#BGEEE\-V/(Hc^)E=(V29\2YYHf@U<CcFb+K>]fFFIf8f/59/4BRA.\53;
]R?\?:ccEL^c+RMR(]SUd6fcW/.TMDV)D;4EFX.8G9#M0^13\Gee_\:TQ2J0BCI0
/(<\7O/G=?-RXE9K/>?,bY@M(UR>=L)#J.LI>I/);=bDR6IRNW1gC4fVc63dXT4+
9>F]1>^U?-HZ5-E79K2#?TaZ]U=:XWcWL-8]#?N9L1V4>]T+VR:b@Z=-53T4.V(.
O0DW<4+-(a,?)I(F,YNC^g1g[WXF&OF5@GJGRSYHOH4b\K5JNO;W[7;<\]B?T5>T
U^#1#Mb+41d2\e>/T_R9&#3L&\A2,GaPKT+;3D02gDfL;(_T6e9(Q3PKVC7,XKZT
O=b^C;P#B&N=dKGTJFQFGF;MC+a4-f<_b/(F45RO9-MUgd+3APD\#4&L;;^4cN/U
5FG<)]+Z8bQ^fWdF4^ed:9>U2#[KVCDbS]YB>(_TJ(JaX0f@/U>/f3Y]@+>)_QPF
TIW(J0E@]>?O74d99?FbbP#b<[<D[S0aOJNA)FgF2M?dRF38-SLDRecFE^))LO?=
1K]=@Z4<GC#;bNB6?DR^SL35bI&:ON+_F,ZM(7<LM>0W6:O_2E-G-YO,8?NISMgV
^.:3B68ZL>-UV6gO^.,MV.0^fF^:X^?Y4<R5S[3PXK#.#g;PQ5F<eZ2__c?[JYNP
/->BXM[]XGO:e\+;0SR^2+f:-403EgH[1dffWZO(FcCHeg(a&1)2bU@K]TUeKe:L
Q)W8c-4J(c(B/E377>2H+G5X7<#N_QS/=NY\/.[[0LP^fZQ:Xd9UfU6Y71#(BK.B
PC6&fB;[>W3;ced_.,Z=^JaC4B0^?24;==<05cd8gAKIAD1]WcE7>KO8Pb)/8539
AHQ[U++=CO.b=GHT5Y1;WZ(#7f@Y.G=]MeIW4c:+KacAX^SFb;8#:cG.[_]KbNAc
8OaT?fKHTeGXY-QJ)(/8I.]U/T#I03K_?d@:)U..4<IFT.O=A.XETFCa^d+?2U7>
-a1?++E1[H<40\UIF4;\GW?S]T]4VY9^ZH.KR]Y9K=3-f]33WB)NB>57GN:g,f/=
RS@)&\KVgTg339SZ3Q]K/dS70gG&8<C-J=BV7]<Tb]4&M<edB<X&O6X4XHK91Qbg
]7F0OAIU?AHc.d:6@GP:7Aa7Q4#?9B0D6#4&fDN-[I=YEW.Y(g4@+ecNY_=Xf:C)
F^b(2[F\HE?X3C/AWK._aHf9YM0<]2#\^D21#SDA5M4(+T0J79=0[]&,H]N\HCSc
L-6Q[YF[PW<QSN6_N;0SbORB5K#]1Cg:<,5X04QI^ZEO9],L,Fe)#ULU1/5[]Tg5
Ue,bc/a7>^\L8F7;M57&e>?WZTVW[)7\G=,>F=RI/fWRbdc?ScS,Mc_B..XUZ#O@
J0OZ\fg3-?(f@W)L_H+[C::,).>9XWHW\.RMZX+NTd])#]=1LLK7dA3-2Ac]XF)2
=3GWGgAJ#\FN;GUQ>5d]a]-^d3O)[BW,4L+MG#4,@5&^-eHV.R(.\.Xae8:eN<BL
e-KZZ/K+::>-XDG5/]cbcY?)2DSQE-adbHE&=<Me_9[QKV<gC,I+?EbJPW2)+D-G
LA_8QP4<QF>ZMB-G_0()USQfc).9.H.+6PTW71&=1[6X36@&U_/T=O?[<:PPX><2
,H?R,g<U^D#c13;8+.D&.:[8WP9?Pf-:/UNLGTMHYa?^/?1OFUI)<?aTTL:035KH
gC>U>\.H(4(R2&@9GAgO:HOX&TE:^1@24DIA;eY5@fF76UH0dg(c0>)f&7_Q2]BC
Y.WPA3>E-2J[dDJS#>:?CcE?64W@43IM38643<?7QZ9NbaJD6;5Of<FMK+J0=Ub2
Ke\4OAV&THgTA&[G\&73WW2-0+360S#97CD+M#-AKfX,Y9=HNSV,6.]Wg2\LC2:K
QaU^+;.C[C8G0JTFM:ZFc&0SZ(baMR3S5<DD7b,758Sg=eeNcSgNM][#ZH)K^?WB
[G>)^=)GS\BCNO2=^U/;e#Kg^eW7(.VF;G[U[;6b,X]T-Z:Te(H(f)4TBEXU:aA7
0(g3?8b(^H4)dga91a:]d^)g/S:W[S]+N7GYE<WJUgN6O?I)GSD\\5=Z]VS4W)?a
1Q\2=IM?+&5_?XM+EQUO_e9#c:5CSJB&IaS]8Af&<0<\9C:+D5H\-fL&g?A?49ND
5TcS4:&7d]CdGZ/?Q:_b][N,8>cF_D1JW2/B3JD\YJ[If1/A82RR9U\;E=DV6VC/
1eBQWJR<aB9fBfQH[aOe/(PgNVECQ,:.]-OGR+10Rd#b#T1aJ6SNYPW?M;OX&X:O
B-DE5^_b](GAU?C/)9AA07#b(=I.<d=7.UVRL3ZXG?_bK8C\@)3#_8^0=7[YK7N0
87caWc-[-ZEZdg9P]Z<f?aD2e)<6?ZS3(a:6.-V&VC,dO\PLgVa8U5dUD2M:RBO;
VJGRJXB_97)@^@&L6;T)I8&B:,5)V4NEFI_b0,3.+cQ#?@@aTB4N_fXSC=c6)IF@
^dcf5cePY_PA<0b+D/6YXCID)b\^Z#2K(201e++V^N)0\fL47VI<L_I&(TWMb\+R
@#EOOJFeaZE&3=Ra/352B#@KJO)4QDW(@J0d(#9Y@1^]\5ART?,=,2@bMfa.7g\/
1;3C3UPBC((FV,fc@RTf54JM1d-dc39H<DG]I_dALSf]HS>W#DK]NNN0=+F;EW_A
YP+5>7?0@R.KF5)3I^L1Gb_9Fd@#YP5AP4NG7)dGNa(6Mg33;L:cIW5][2[:WK[Z
+L,G8dS?DH]1WWBJZ1bXfe3O3E^MaeZ>\@5_#7X&^3fT?6J.CSV\[=f]?BgR6>W5
(gHJO^d6)E594D,#;EQd(Dd+]3648bN/M#5J3;&_d+PcV6IBCRN[@S02bO&.J0U1
\B/.Y:YM(RLE6CT1Se5:/_R:Pg/e[aPH:F:MSJ46425G].?DY/W\69ERR;+-++=d
aV]-^Y-DU&05[-QeU??UY;<gKC-Na2fZAXS>8JV,59UIK;>Kg0>eV2@>\,]eJ]W_
T,@,S(LQC)OJI0d/=aN7,5cGG+><O;.6Xg2d9ed34dK,EaIVd^EC&9g0FOdHUT1H
(f4^DCHcZ,9c,eXXa8Y:aLF^PP\\M7<-XVdNC)GB)U:I8JVEFY5S-DIIIfG2/ggE
BbOL,2:WKWLF4g(I,[=6#K5EU3\I;#W1PQ_&DI8d0)B:E;.Y<-(G-)Q63.5_.=F@
f:D)@K+[g^WOFMS\&(8ag/]@V2d/#<T5AR6F;6JE+-JfVgUSI(+GIL-/\<c280M2
]#LaZJ7KUICReJfece=f:GMF0KH]@a<)[I^:ZV\/KJ;4U7NR9fC2JV:-=L=,9CIV
1M86cbC)R0RCEAC<d?f7(&V;CV;(1S64VH0+(c<6^g48<D.X@J.6Q[3#N>>:)=DR
[QdTDBJ20DfY]8VT1EJ.Xa8/I_ZMR;Kd5M),b_LU20/..HY^)dcP;6[]@0fNV];F
EII#T:S-HdXC.QI^O&>DXPfKNAQ?Y=25Q3c/SLG]f;gK49H1KLN(=BU.[RSggT=8
-7TE8<D60.Y;,f+eI+87d4?Q5e=9076A1WBD\/3<Bf5CYSRb=3MHdg7T5T>;:AP#
fE-Ug/QM<PbD(\dbM3:<DP=9\5B0?)W(RUV57Z;DQRCL4M9^.9Q<HP[I]0ba7A(?
0O:>409GL,YW>S=16_;61Pc2TB5?gDDJ[X@S?PDK//;WV9&88RcU4Za&CMF4VH69
_^b2^ULPGE&<e1_7#DOQf?I>HMae+AMc9e=9Z=TQV8K5ME]TCZ1MKX1VDYC5)=Hg
a4(PUK=/\K=1Ye1-+[EL2_-ZcX72#W<;bb4<dS;M(;LG^P\LQI,-@Q,YDN:>0-1.
;EX4W1/MYS=)V..#PX@MAUd:;5A4MIHT8@KY[F;WIQLM-#b)Y,GEe9MPgDM7BTKd
<W&:_AMcgOe9(&D\R:0KOfbSDU4)^?DELF@-#TdIU=.C6O9WW9XEa:Q5O8[If[?c
).&3QVNXL.U<M2[6/Zef_&2dZ(<8#,JHB>EN5g\KHHWL9Da;FZ1JF50.XV;IbPZW
e]Y6@YA:E3RI^+Qcb<cX8ZRH9?g>=BKR7[WB6.d[KSg@fXO&8bb[H#6UD5DQRXC=
H7X403Z:fB1a=OF\3ZRU@#fU8+YR[YT^gbLAX/C7[PY[_/C>b5H2(\a&)=<4I<EE
IZ?\gA(BZFEP3;d[Ia&<QGO_2).(W(LPdQQG^g=DgP/UeX2^;E./3;#E_60b35.-
;/VMHgb@KYWB;14@+5PUE>GgE-g+E)5aS^.,fQA1P#N)T]MQ/]4=3(+]9ZDacM,<
YTe=^A4OT1@6M@=3,^Q]3QUJB5gGD:D,YC?(3_9/8W:_XFEQ2[OKOXH.=ZVU#JO?
aV@Q@-A]^7Q#@f#Xe.R[4MZX+^3?g>[<90@R<BOP=<:Sf^N8ZYf5H^gB]6dS6dMD
(b..IQ8VW3-(Kf7M\BJOe0b#TP8g/Sfef:R-3K^JMO3=LWDDggZ@68I)HcU2OE;d
FDLc8V3EFPOU/1Ka):44Nc1c27)/d3eS^KD:3CL3dT^gJNN/KKW.GOM47FF?/C8\
\e(ASMKfg-V31E5;JL.\0ZE3IV^X\6H2Q9II=_I7B-7FHBUB5W7_QY98BB3JBfT>
cDSU4-&+B8_FM=VGA-)=S#dQMIb4VM&@)>)S@+2_1-UY6N^-+N\UQ9@Y:506I+.1
0__(dR>K<^0UT8[1297@@.AWNe>^De9H>cb,Z5d9Ya,KU5NRY-7bXEC-XFfdC4XV
ZND).V7<g5S>RN?W&7#1=4Qf2OZfNHK#Z7(c=@KF]_@f_c5g4/]TLTeReOfMVS<2
_C7.=5R:b62VW^?NP+KAd.L(V_//1_WA<\NHRXeL1I9K;V[:4bf<eUB,;S-GK7\\
32XVKVXJFI_UBL>A4a\b>5_0G9^H)DV@AU-_6Z;YM6]NN)KR?TYT)P[P[WP6.:c=
6=>)]5C;=L=dWdb8MV.^[ff=O1P:_1WW9RLIb-cRUf3II(\:TK-DaWG1;_dP4f5G
#FFZX<]H@IEa,CL/16LdLG4BW;62b@P=g/H\RD.#]4Xe78YHD?45e#UN<_3\g[]3
X8eVgXN025OaQFI8-,G6T2(bOG/PUA9175\_OBd;a/E/DMJ3O-;>ID>EM#>8LFS3
?=M-S.,eY8NS\aGaP1gbLJ:=2=f)c:DVIe.f5GUcCE#EJR1[?[RLY<de^LJ./5(@
OE&^QIg]3]<RV[F-<]H@@#58+LT13H31T@7T-9T]N^FJ;8IX(,ZQA&]d#8+ZG,]1
P3F3YVJMST@POG#G1A,2YfN#7fIVB<[a7I[Y>AN1#0NgLWc1EI]fS6f0/8fP@SeK
;C_+-[(/(g51Be(.4G:T14BZFHE&>c<S213BMf9Wg0TAILTY=RYHN11E)dRMDZ\V
T@H)?_A\QCF=LLUGaJVTaDW7B0-OeJO/WWf1OB\T89?WF=LWSTdgS:DR?1OH]&AT
G@f22e^T(I.e-X=IH;^,#>,M5Y4YJWQ+16TDQfDH6<ND3E1?f;)d]EKaR6(X1@E7
ZK4G+>87T#4HY^ecZ2Q=O4G=8/PcUKYT9W<g,[X-\CI9P=O3-b)U6WIA3Z]5_Q[6
;XUaX>T>:=E=_g_@T@(CLgP7WU\T5E96@-KUVC_[d^?cf6U6/HdILR+6Z?c1BC.\
THU(]UT\/Xd&H9eMI<_J^H3QUC&B4I^1<PVMDZ5(RGEUUB3R/75;<K\aNVSB61>^
U)7=4F-7Jb#IZ#36#Q]gJY(-TZ[)L5;^dN3/01WVAKXD9M\9@QOe[,&/3X/0KXJM
DWfMW2+c-^34VB21aP[>9ZDO3R)\6US3(1&a-OgRDR79B+SL+5[EaKW6_Y6U6F6d
a8gDMSUNIDO(]&=d+U2&8D85U(J-MH:;F>WDdSJ&7f;K6E0NLZ>dg4PB4HZ5[dJT
K:GT&\EZQe4cXU+Z?O]9McVIUL7(E^R3R<HN@]MDgYJd591QH[M-(._)0.8;D-3.
VPbf/V[<,ZYNf&:La7@]CTX>B+_8P2OaE0N@<Zb&<R96IVd-7V<b[ERS1_P[9.]e
??K=P8#WN?3?e?,LBZDLeN/MBGMCeVM4_7_5<>/;_HfF3Y>>#-K6#K7KNA[VeGKQ
M,7A[@0HUU>3gQ]:(37C.PCZX7>G6TD:ZFC6.;f+COJP-Ad+g3P(#LZ(NLORY_-G
FK#3CL>:e@/3&,W<1K_\,X/:>SM:]=+d_G9dYX2VP;W\Z]9]aETCG&67)[\a[d5X
>I#E73[bPe2FLB&>:@(123+B;f6IeKHWBQQS&+NA/[dPIX(W8QGDdVZ)R_gECCff
[aK=.^(b<2(LH,>OJ#[3Z[>L^(Y0>G_]c+2dM\G+QKFd/^<@TQ91?TXgI5PeN93Z
GSI>TV-3D+-Z9e3RCV\O.6g6YBGG6D7#gb-b+V?J4DXTEf;,F3J6+[.+J?61A,?/
^+(SAT.Y)A53<?d/@,bP,M5d2,,LQb<;bYfFf2&7VR2<B\C1C:a/NgO]gY4;Ra)a
OVI3/_\J@_5<0XHJKC[WO76/;VC\3a\bK29G7-J,HTVNT1-J+NYBGU)@V-Pe]HFf
@WSWMTK7Mdg#.bJ8^d,I4QSDec-E3I0#G?#Ua<MKgA[=VFfUDHI(87gf5;e28cRZ
Pf0UfKeB(K4XQ=8:(#=Z5-2](XO/d0J(c<JbBAga:#(IdRS9C?G;=:@YaCbA_4VO
,HN6-T?0=I#K<-]HfL867SG:.@Xg2L,dNLQ:fTY_V)6gMK#UY\\^Y6/L@a\2b:^4
L:a86bZ^\U,G;I;BS@A;-ISI9H7bR\XXP;;Rf34,KF&1K:W7QLU1D(TH7?<BI)cW
WU[ge[1B<e:ZB8.4Rc-a&#+eCOJR=Q+^?(K>PfKC^F32I_dOE5]FU#0IQ[(;b/<>
)QZP<J#0dg5/4JQ5H58S8JHK-Q[DXP]Q&S//3P>9]ESU9YWZQ@d0G:Oc0E&@3>IW
IW?2If4P-\C[O4[XA[JDXEfbNWV#]]K=O+Y7@_/N&L-F?AFcQUIE?VV4.WZ_XM#c
(.[]c/_(E?DX)<LKST_a:S2/ESJg>3D#?f(^)L)M2f\_4fJ9-Y.GM]7ef8(S9Y.S
JM/)/H3A-6f:FQ.dQ5e^)bWLJHL&c[TGfEE),=SBQ?C,OXbg[7B>S(g/74gSLObf
#:A<@NJf;#d&6)]C=M/;ZVbRXC^03K8Ea8ea3<GOa@FZKU]/791=4c+?5N9U)0UQ
.HD.]d,d5V)0QO+9OJQK<R5&-fb7,:^IP5HPB^ZUH6#3GG;(@IN;&P>c=10,0+P-
.NP2>)72J^D#_>1Gb0;T0TE+84F7e2K=ebFL=bc:R(M/P8\=T-Af\ZKW(XB>C^5#
W=7IQ-bF^e/F(QTG:OZf3.I?G1^&30C<B)B7YCJ5G5]gWgKb;(g4gLJ=:7X0Q49T
(d.UePP@[/O+,3U#;OD(Y2^Q?bFg21=35DAO.ZB)CUb1R6fF04)&LP+)_<7NE62d
S?K-D^B)LgLY)P2fWB^V\e:R&c-2fK]HQ6Ha@]Kc?NJO))L@ZV3GQ8g(@R2YCacb
;AK(2E/EL=]ZWA\OaTe\;\0Z.(JFIN7+7@91;MN8&L\#/b)b=SabQ.FV^fg<QcDO
.;[MN:N9]VL)KK<:F0MYb-2daW2)7/\+;[+URAgc87fG-2@@B:2@MXXA)-a^[AH_
5SG?MTO=6MZ2#_?.#Vb8^.F@:a05<[[4<cdcUR7\U7^WJGCPN8U(0?LP>\1gI^fY
5Z1GYR_A,QA1_a[9-fBNCDV.eH3a,40T&];WcXU7b\bS-7cQ(cI]?O?ZDV>Z.@Z-
1bSCZGCJb42dV>:((fOE1^64Kg0L(+C-=62O+4R_#K-9O?H9YgZ[Q[BPD=d065F7
@G,]b4I1XSa7KB@\9MI@WA)X.=aX8FUe<6Z-gA15JLO+-a@HO\aJSO?&aYBCL,aB
U=B851-F2;N\\;L3\#97D4a4^LW23gADI0[cE6Wfe2F<EcR)+EW,F)]R@KX<ILT&
Ug:3J2AH\7H0G]G>(PbLQWQ;/E+K,gD;39e1?W2KD68?-U:#<e)fM8^:>7L@#fd]
DNbU9..^;Cc0>A@STP567,U.;MH#+bCdB_FR7HYMZ(2?;fS^T0(4)[9g9)2SX21>
LA\;/D+;G.c0?M7a+LT=(ZD^EGFaQJ@6&QOR<R2g#RMO@Gbg^#3@X)eIUL^g\C=/
>GDMaWC+d(R60VgcFC.-:Z@:bIfK0Q\\_NAZN<Q&3&8e0:Z<+R9<38-IdVK5c\H>
S:).4]9/Ee-ZU^eZ=^Q:_A7X2IDHR53HI88/Q91>Y_PNP+\DJaMaA0K<=f0=NVPV
c1[7UGf1d_VBgF89Q(N9QC\V[92[c_5@K]DZA]f=NK97UDZ+&)5>b.4_?GfLCWY&
\4ZgGDHTGEDNVbKg#1Z(B##9_&6AK.PK1aaB@W##caX^?Nd3J\7A_a.d<b-1@eF7
K?S:U[5I[&HE<Y5b(Zb&-AEEeZH4]Q-:FY[T^J99L)UE[7/M7aF^W)aU4[8Y9T[E
1efVfL@b5T,G\6@KNUWVCO^Q[cUS+3]P[,[EL#H<2Wb84&1MJG^T(O(1NcH3DTM5
&B9OIP>PdV#L:I@DFc8cZ/<8^G6^GNPEQ:H,0X?Jdc)f2^>?\7cdQ+(O.&<??FcX
]35SEN926Gfc)&>NMTAc;LbC/bH;^PYe-\@(M3.f=G?P\1=BSTRIOOHNg<1aMW^?
@V8d\<ZV=72Gc4K#e/=NeQ>;=LP^:S0E[+;d=/K0>3\/^V42151NICS7ecN+[@[C
>-<]O0EX7E[_g1L(Yb.:<cTY>S_=S@DII8=16A<2.[9N,E&C9HB[2\g64;TJ](b4
EaXJ_<<0P_KQPO<89:75Z3@_YV.1:QLF^C5==O-=_Kf6f^G[8K#X=<U)J(1_[V;6
KUQ\/eARCB6Rd-9c,=\KNQXJ4SA75VQYJ&EVaaT&f#=<.(7b2;L+ZKB.<bUB^f#F
_F^K[L558B9dJ]ba<V6/f<cJQaH@610b#UN-AMPP:T:?dPe+gVU\ZJ;21OABCS5Z
FWC)2WW=[(g];2MS+QV4@SVPPcIH(B#^XMB(<&]HI:?_Wf_DU@1P@bMZF#XSAFP2
f]b^J[C^eCONC-bUeddFFK](J>K5AFW^_A=2aI(ZHa<4^^=;7M;]U2,g3KL/>+M>
>A+^XB@/Mf=6&D6S09=g2G5@ePM#++:9cRM2_]&WMQeZH02TG2G<66\Q^^&XTa_W
c#&1MfAR+\>dB,C9<f(JM6BI8QAcA:2?.XW7bAP/_)aaR>32.E2=MaI5^VV;4Xd+
NPc7;&(G@-@1]#(g5Me]SSHWDO5<>+D)R1#OA[NfTBe/9LR<f?8/08aK(_I12REJ
JDaW#NH4&aU@X3dbC<:9M:fb/E(BQGH+)>Y]HR#eg8A-E=-WJ)1GVXcSS_R/TTc;
2(#@]T55JOQR,&JA2b?g\<1AV[MOc/YB2aXI-E_YGWZ,We+[;ML7/HY:#DM9UM)^
GY:Zf1@g7C@S+/0M@>Q9#0g4-6),d&Z/R.\5<I2TK3CUA)MOPN](-VJ1>;-2L;=Y
B;\V+8_;b._W@=376T\-::85<MR>OX/?/7T+3?<ea[a6LLCQDdR7W@2c_CeVd<VB
](,HXNR>?^-,e&[KON4]6e4TACIYA@]3GAQ;Gcb=CVYgc<YA755P4I[9=:VBf3Ea
RK5+L6K7Y\WZLXXecTbGJ-@;bf)9OA]B]4:MV_3(27J/DI+HZ#\<,0Q<)Ib#M#\=
<.F&(0ZagB@<P^?5\Le4PSWJ-R9Oe,N)IH=H?d.KLCX1V5.V(#U/d^dP4+>e2Y\g
(T4NM(Y&.VDIV,RTa3.6E56GF[S\L>R<f>_7ZR>OFAaABdE5PC+#a@FYL(XWE37e
+]#US#]@T7bP-a_:6/T<1#]Q2=a90PM4g\/KA<O-2:+94d^3<W_?W@+8b]]d&N]:
NLI(7K0e163AgH.XC)afE?Y_aEgGEg^K=Bb\9RcIV[URF/c@De.P>3FT?#2Y;O1<
0_[ZV>DEJ>J,9S9]L_?(g2aKd.6_O\.ff,T+B@.C?CQ6.PZ6^A1\WWgQ^0;RNJWb
L&UU70aa6\@-6;/3:=I;T<:@PW7R3]g8a\;SU?Ge-#>3,XbW8,>df@&[],#aACC?
,cP<CQIa9/YK=[JcML;+eW>_+T-E;:RQI]PIEGab2JBF,Q&4gO>aX84_(P>_HOTX
7S1[+QE,J2]-M/O;IJ]^U6;FN9V\b/YK3ZQ)6+U6)][5SE_JO^\5(+0QT?G@W7&J
cBTJ>DD^Q,1V\?e@XQdM=L,T&E=;(.bS7-YWe1(FXN5XHdHUgWJVcA:c:@/S<80_
X_MO?&CJF[>?+0T+5f-_aCB4fS<+E?U_7\I6P5T_58NIb8H?ULWI9,U55gNa44Ab
,aR5f(VUDBC+ZQ+fXPdeJBg?)ZW@:a-10VRM<EV&J5339631g<a\JL4H3>X+eJK5
X#,2?35<)^\d2E5M4.Vg/&Ba1WRFdZ(?UZ4Ge12,Ma;U5A5T.Z+ENE;ZgJ@dPf/@
(8:4Z-(+\SM2ULDMb#A>(NP;FBKW[)LK<(8+EN=]Z;2@eWU\d=b1.B3ZfV=5B,39
)gA7^W7Oa[JHGGK-52<5-JQ)5BbAQZFcM-6X+\LEBPB#C0XBU2]R?cA.FJXb3-KQ
9PdBgOPI[WgG>>G^Q,O;]WJ-)HfF=1eO\AB46=XEMfXFZTJQ39W4cK2]LDES,O.:
#C/#eWQK2A[E_6,SN>RJ@fS5KPD/Ng]_J)X]WONW[^TJ,N^=Sb8KaN^d2=Ia[#[T
f]Af,LKK#bH3+\=MdU]VN68MJJ[Pc\\6/BccI,K?V,19;E8b2Q@He\E\GW97PGIS
.G8X-g\fWP68H/U:79af]g]O<MMY[[>DbYL)D14?UI6A;WBPOG:eWdZ59\?@)0SP
,L@0.4?I/TIYdI8#QDOg#BfUVNFZ@Sb(TKI2I9M17UfGL?e#LDIa+=&#+Q-/G&Z_
NedGeF2^dc==QKc1S+WG&ICM#S/g+?=<SOGULQ=M0GC^ONWZ55g,UAPKZG]9?XH_
89P6dC?L(>IRHFV379UeZN)PAA1ZJ[W_H?Z5Q1@)IE<c8@_LM2^AU?9ZL243?cHB
JDRKB\f8HdMC#0;QfE+.[A,:bHAJ,0,g)&?49G4KZHF>1L;OS@73V3=0SRFO-]Kc
F4MN<ES2@6efbE7N,Cf]c]-JeUfK8(#f?X^@cY[L4aEWGFS@&?SY^K;0-N#0OU_7
Jb\TW5-4LcN29JIR#=T]]R>B(YVLU/ZP6A5@\_=5<>AfB1Q6fE4_fAF8:?M6,Pd\
IaX2MZDH9FC??Xc_RcOgD8S]gUZD40WX++?CN:41#-I7XYV.W=VdW#FaLYfLQdX)
[[W)f)N:R:5Ue]ZTdbX_d?P0]TQNNN.#H_U4X1<M)[AQCU+#A7UV-2>^V#L=:K2#
WO7\(?]YJ4/&EAg;7(PS+5,)[()#;:@-8QX85V?2_]G8H88&-e_O?H4<)aV\\-4T
Z80IU+<>;\D3dZ,)F/5QZYg8;AfI5aJ(1dJ00?/K_Xd@f9PR+QG,+b,BOBM)2W-C
.#XRZHb_4>NWUg5eYa9>NU7&EP:K3[]Y+3=Y#Pc2IG]OaJ.[\UT0.<[f+b)O/H_-
d7(R3[H5DPJTcU.TD4)CXH?6Q8F5f:20MER89RT<EdJf/@.WOFe1)GaD?AAD:W=E
Q98R-9J?8<71-#,;[]Q>&-3A1?e4[1_GLdP&1cMY:>83fYa#\Z,:,#QO;&_PE5/a
/GM3(UC=AW;>Y[6eD9>Y+g>GRFG4DbS64WC8gDM4X+UN8WDg<A(@DR7TLZ;.HMLZ
C>F0+C>-1<W^0bQYfcWfA.KEG@FE[6,a4T.0YA=?<::SK@,3b#4f?/6]<5FHF8,]
1-9#ba_[Cb0@8^2=/Y?/SgETWe;Y3V&K1aUCagdV@gYY5L)c>U;^dDYc2QXUMg(,
;MNJOC?>^4RA?],^3_\[<TdRR7B3XDU&Fb>]c)R/RXQ3\\0a?6<WKWL:COU:I#9:
S8YaO2))\-L:T<ZT,;e,4LN>FBI>gYGFGXH0?0CDJH6]gCJIaDd-Y_>BaO#&5+A=
(Q^]Ve?])/J.\gZLSf&1]g-DcF6QAf,\@CQ3OD7XG-1;fUAI0I+953SH0Ye50#e9
P8CZ\[W.ERSeWUA4OF]4C7_[S+;+gQN<b@[3,0GZ.-eLC7JZ>ZV,geO>bM^]Zc>U
Jf9V@EUQ:7)]4/JaQ]HJRI+^JSPe(UV>Bd&W9YK6C?M6Z[/7dZYgLaUIXCL.76>F
297:QCdZ,V:6T=W]A78@=.cVfS0LZ-R>V9OcTWL3JCP=JS-K^QR=Z=BNgFDKf1=,
CG6cPAFT.[\:/)GOCL<4?KFSbLG1)A1IPRdKP-V=4daY[5J>/[=RR10>-&=V)@2H
]aVXd[7XbW&W?2T?WbU587Ia1P@0Y8;K+BDd@XZ(C=)JNBBA:RT1]Q@Pa:J?Y]AE
<J(d_M1M2N>;><X2\I1KU;[T@cYHgN/?G).:2+e0TQ(8OeNDGM2?4CU-Jg]b=PSI
@8>QYGe]RM_UFA(A87_XXJ<a\[_+M;SRP_FN][:IK1DFQ=+XfV9_#:5Z<;>])8TU
_PgEH@:+d?<5K-V;aV=(1cb_82Xaaf6T\UMdNS8e.>2F^c[0HY52B&.7J5OGfIH2
K:X5>\:DG\Z,2&#HI:ZOfUI1]R=EE9?8+05F6BQ@H_D<5cedMbUNHfA1\_9S:D+J
NH)9KQH-db96T2U_e/5aa/&TUC6]YADYfPU1X6bd#?=N_Jda:aL-):H6^gRF<M</
eQY/9K^=L4N4[1&&ET^YWJ/#>UC1PXX]aCJ:N(&&?7)?Ife)QPY@2FH@25_DAE:b
&DQ3VG>Z&)/X)NfOfB@+.5QJ\)>31Fe\E9Tbe)W\W22)[_M:)/4(=YJG6.2NcO:H
XV^<ZPJ?fIEF--Fb>^?B7f54LMf(dZV;YIZQ^FMc0K95F^>]gYP0,c\?_U+OJN)T
#0DIA>P[-UKOCaOZ^P.1Oc7H@)GUG5I=FCU/QMWa<ZUD6gQR50d4T-dKM(Sf+0d2
1gVI(KXId,,\>&7Q8I2_R/dM<[O7;)O9&I@P&8WS=.]bVY?1Ld42,e_=+W>_VbP(
6]S02f)-DZQ?DW_[9Ta-5:7P4=C2-WCQ.M0eZR@:.:24deXRb/)\gJ;;7,]E.=I+
E&9>T8H6Y-US;dLR]@/CR:f0_\Oca5^=IZO=P)_Gc.H^DXcOY#>2YY^SS]@<N[S#
6=4SC(AH7d;4-A.][CeMOY]Q;G7_G=G9>=Icd=178>;8Wf(a#GVY:L,6Xc9JH^D4
(fAg5J_cdZ6KSNYHOGc^JXWTE=]bYG6ccFf9aJbT8>_X6,d<P\EW+aIRePQ3YYe;
c\Z\M7JMAI\T@cV@:c9PPT5;1RY2_)0+F?DX<;JV1KFLdO;QRJ)6b7V+(H5&X;6,
.Q=DPZLNEZ)H+U&EU1HW]dF,U^ODDJ04FKU+U.#OT7B501BZC=N,Oe;SGB1[6DH1
c;>FAQ/c]=TRb\YSG^#N)^)IWB]KC8.D/XFZUd>/U154,VUT4\XX0/M[\R_@(U\C
A8Pg+VaV;(LVAPFa&ffMCE;74F+TdK3HBCZHC>]&#NL4-JGF(KZO;7.WO3KcF(HM
RMJUcU:@deV7?HD1S2IEb51W>BU/7E02YHNH6(#>+cI5CW@SMKDI;R@:\+L+C7L)
=a^0A4EgK5[We.4aM,GJ&@L:CKZ,,\#00/4^(NEfdM,NSR@IT?&-\H&-]CKdG>\c
X=]9<ZEe,g)U.\B.Ke<&3NVO7c83#2SFLg^M0ed?26a&.,(UTST5P6;5PAQPSOY3
[)K:&Qdd^JAd_^NaaG-_5FLBS1=7)R/AY@TDMbcaNY:RCJDJ((3[_^0M4UCG:]:c
MNWI;X_>WF;YQV.)0AW,VE<&XQOJP+=)VYI>7b+C807:HNdXTd@8]5EVHY<aKU3g
cODHV:<IA[4I[]S#OJ-Y&N&?/XI7;Pe<PMA4TLQ<R_@\ba?Ie2DEd#I#W(1QUV2W
cbS,28OJO.C-DH>L.#)J^,5][\FR/5)F]0GQG)VSGN^X8SG&?N[R1A&PAJ5EVRXW
:CZ=<YR@RF@Y]-#?9cEY/cGfdB9#C/[V_^@3^MI#,K-b8@eVOg#M7Hb6,\&dbaWD
PD:M+^dBdg65,>R-)^F&PICMJ91#E9_)(>NMO<Ug5bA\4_M\<?3fe(LC6-EBdP#3
UL16gN40Y5OYIP?bSeb+(dg6\be=UOW2N1Q&<2^Q]0/-NZWK_#afBL;D&e+gFU7A
CYcbTfEEX#?9NPH9O8[+.@\?L?a:751-VHc6O^c#QY7IVN1(3.FW3cF3JDGPJ=Vc
4E#1KMZKf.d3GIH6?>=0BM>@.RgM0&X/)/?XB/DSgHW9I4VMcJ4X_H3AY=QF6L/^
99I,.X4<Q,7183-U@,UdE&J2,\&_>Id3@KP8D>A+9XE6De-UZH]4/Xb7eJA1f.8I
YIVHIg2-34VXPgU]FbBbLF;CX?@:/);B@WHZ&N<;<T(,XT\eZXZ@L53G8P(-[ZD@
(g_E,9\M1N/Q[O[I,1&fX-B^3=MF0b)cL_BHO;)@HRaB8MVg2#I[@CZBK9IPV0c^
[Gbg1Q]abccR5dZc@3<AU+=R;&_II]2RW3I_-MA_B<))/4:&(MQAXeIF?;fMH+8M
#X:Ng7_^_dL&1e5>gXK_dE1AU92K5WD/.];JYH#FGY?@g:Xf=]RKJD3d8dC[7a/?
4fK,g(LR2S&O[&Hf,KDV5Q.R<2SdI?\)bZ58#Z=Ad6[<M)R&?)I[UcCOgd>Y3R30
<1W]NSTJe7?):de@fe+UZc[gSOA#c#Z6AgX(UX2N9#NB=eX[]aK,Hfa5KfT:VR<X
2<U0QG#-UQ:8[NDJcK-a5gVL7YH:aF.@QKc-]R?WY3)0]5\<>SAXg#1>)JB46f.P
eC]?C4Q5gU34Y\\(2/7P2,=[ALZVV9/-.JC5DC4EeV3RF#H?K=#8<dFP)(D:9f;K
Fg#D-C[PM?#H;UK0#g_)(&WAO<_R6d]3TH2]7,30<d1.g(XabD3N#bL=g[gZS72R
/TWQL7P<(4C=)7:<@F32\Y,\01@58<c@M^9K,XbD_N=)B6WTO1_IYff?&d<_JC;9
1U6<HG_&@:dFJ=&(#Ec,C(&C)3R\LH?=?EV4f?P\#+ZK)SQ#6c/M\UC>@Hc_/ga9
f3DE4O#_6cfTK?6C8Kfe;W3DE(D]&A2[XW+CT))8;-T:1X4ELEHIZ;@?,PG.8d>?
B6YaKFNE3eFeXa4@R9XHdYbc&_45dY:Q_>\9+ZTIYAf#A8HPDT@RbFed^;;+.=NE
>?Kb<2\M6_B5Xg.4^/8[dPbdSDL1J:D.S<0SQ8&g5]6[Q6#e&]9d?Ge1(7S?]a\5
__N-fce:NcT>O^QU1g@Z5ONZTdQ:1W1MRJA^A>3Q:1?QU))X9BC,aFW<]Cf=)+CU
GML]fWTcdUL[,V-Ld=a^:69N7@B;\Cf]@N+dWPT^a[][IR(;O)2,O]Ha317L](6(
R6RH<ddeAX95[[d7<C)1bdTWW2QHXFIAJ,0@#ReH.K/:[)-N-FdZ/B#^OEB8bQES
3]-V3QXLQ+6>-GRQG,?6bH8a_?\c3#2&fbP/gGM2?g9.J54M^@[76fe^W0-08M8<
O.)\@(X<[VN)[aFN7-LN]?J2Dd&H,Z1K;4U[N)=T5O@g;GCO,4gfOGX8?af1PJB2
(,L<g-Pe(TXFJ-=Je#f7WaeaWSC.9??#:;X+bg\MgSV=[IYF0+?CQ1Se?\-3;(7F
KJV_M\W?_\TMJE/CN5W)@AG&+?2M<CFS:IKOQI1Y6,N0KFaC9KgY]W(GUF7gOUK0
OAS5S^ROI).aB/G9N&5^:(,JHCf[DVJbTK7^,QdH;SD.f5g1aDY\:/,Dd;I,]LK0
CZO>dZf74H;Q[fKgT4;U21H^QAZg2CA55,NUVa3.TZ:P#1H2W=-SALOPF>8[VQJ]
/f4#+6a4JH]Q#IB>g4YUO:40L-,9]g^?#=&;DLeR_,5ReGe^=_M8c9[a^=HESSW-
?F0,aH3_ISIXDEYZ2E+Z5LZHe^ec(W(]@-AM2-=C5)WdCd<>V7WYXbfH&IOTZ:VM
E493QCA5b:BbTFQI-c^QUQXBY[#=_1-E#CED-N/7>?1C>678@,R<g0:D3>U?^[/[
MLcYT@2U\^&J:/0Y92VVJaQX4Q_.1B0M\VXXHLc\D<W_f^^K+@6g79NW(&.2QW-]
UVY[NG@1g(5<S89f^X0B2W)^b(dYJ+DG4-/0B)f/^A[.[7cT53.C(7;A0T.4/KZW
T_16X50/e#O1N7(#X75?Z;<2fI#[=?6:fUH,#59DRYFPQ@72B)eT,bNW]\J,M]/W
eXZDC:Q=K[YgV@d:R?-)]8U^NYVT#f94N4_I4<MFUH4<:;POf-:E[@I0=KTAN;,Z
1&#>-)V.CASGGDcFB-J[,?N6O3^,(g.JZ[1]cX,Fc30H(5eOUC2B=[W[+NHW=EPD
8;ZZRg/:>YR&/&IEUEBM#[,:\8;=7&f(S5bM8I_Q8JTXCYJPB&+:/A2&+Fg\7-&7
K1M=O,;=FJX>ReMfB6W@S=,gQO^2#.YG[e@DREM/g@0)a?KD\f;YESAW^T7R9>fK
NHJC6US>(KeS_ZfA+=RZYg6IK<G53g_6#:e6cV(9Sde_/KW#J515,-9XEFE41@UJ
:f+0DEL><-/[[,g)F0K=G>G)I#e^gU,_XTb]UN-gM/OEU<Zb/FYfA?Oe-8+1QW@&
T8I]\-18DR[4IG?><40QEAgLQ:[bT1D+J/_<32NPTH6^<g@1><)):Q)[WYAD/c18
IUAZ7;WU<M(6T14a)-J3>WdWQ#>f[c(]/e.[XUa+0BN[Y<eWQ<f6b<J5cG)@aRKJ
6^Gf/,\SYQ3/-[3(Q[J#Vf4Fc][OEb1Jc;T)_K(36Y8Y<G2:9a=b^\:JW&gZdB,_
&8DS8GeE)#>f7aNP&K5:T<K4V+CV@&MOTWaW0/3@-IbA5QZ\DOFg972,\D5PZ#^,
D42C3\R#RcP9?N5;.,9a7P8_VD(:d=7H/=>2])a=)D:5(M/FUXMLVL58KBU[2R]7
-Hc?J7(S+Y:-Xg,8BcE2:c5GMe+#,^_?A.</0180Z7@OYV(.4G3bG?2Sa_?#C5\C
B0YB6TTB/(UMcdSdeI0fD\4MgT/<AY2>-f3:,_<X>1B2S(SODY-@?WG3CZCB#5^f
d.-^M_@\IfL0T37TP_a162CgQKX,X,2FT+d/&U5JP?<I&?-&QdBg4SZ9#0W<,>JF
Va7]cY-AD?\-]Q0@b[_H#R1^=N[gcK6YL&TG73W?dCZ2EX<&ZdQSIO0XZMH,7c],
b(c>g.Z3DW9fg;:0:17A16^5ADZ+-:91U9eLXR9,[(>Q<)@XVII@FMPgFPUUUI6I
XKg8OK#-E)L@[</JJ+A(ZSYU0.Y/)3\=26[P.^94F2W43c8MB85&4XV?FZS.GU9Y
)PBBde4Fd[)B#BcBE30fff;8>VJ1K&))3=UgIa/3L<D])P236X1<?EO4L_N42FG7
-3@JCRQU><g#CQTKWcU.,/VLZ/1eM(IL2e):@_<8YLG8(0:=,R[H9RL#;:&Zc3VT
:FOWbgDAC;K\8J>Re<a4<LW)XN6c;WI]\IOY^Z[Id1(IKdMD&(:3G/O#bKd=Ab79
>Eef;CJXLTM]7.=GBMHFZ-A&&I5IF7M88FV>(#NA+C7.L>JUW\B9cUV?f[+.D;F+
C_eQgNQ+8^7EV1<1C.Z+Q@gX)(#E.HC[bdTG#a-VFWLKPfW-)RgOR7],]ZY<>H:E
Fb):NVBceS99I=YPf;685_N0#a/W:EMEQ(d>MWQa/-NS8X851@J)OJB)P;7..)Z?
=b2KCR7(OQ.LJ/73[R((K-,,8Ece)8D83T;DSQWY(g=VJd??X40:;H.G=8bP]J,+
X/;:7Pf,/e<7+&g<aJOD7dZ530U?4XA=RAK3<[(+OEI?cZLOVO2>W;]TN/4U^8g/
//NL0IfO4Q.G\E^,Z::-Uc#.AadI9R3B.H208)/a9KJ8cc:Wg3]LdXSH]Y<K?>W^
8GF;MS1f;)SEK6XN9W&L(3.@aH3WW?WJaKA_Z<g+5B).;[B/-MaUAN_&egDIc\B&
AeEEEb;=0+OW?C4KS+FVV1fg6+2>,#0]EDY?dE+(2Rc>U:H1X(K@3fWfJV.6J8U:
:,K)PR#+WF9/dP40\)RMCV1O.E+R8H\b8H<+;BB]^)0NcMNeR5-H,>6,[2VXB&6a
K.DdS+&XT?Z]OBdIR)57BAcM+d,F976YScZ=J83HFKO&6[O4;VVb=QgS8?#=+BGg
B,6E\,B.9]>Y-X5#e7.[MF9Sf@DDg/7Tg9J82I(.&B0^5BKRU^PXC,dE@9KPJdJD
@<.V=F7,Gg-V\YZN\aW^QJTQ0_/E#9XA#4UF.[0W=>AfJL_H0V0/RH?_/#>RC7GN
30J-W#DdP6?OTMV2W>:b::A>-;QFV8&K#YN;/b1b3>AK]\#KH=J1,#VB[DS,,QN-
0O5gL]ID)ON]fV1]Te\SDR+)V:9TB(_?@&-LN#^ONeK&V&B5Oe/;ETQH2L:Z?CRQ
V\_Mb1510IAd[e&O>SPA1ae)UK:=],=[_fKc=6Ha\aO=;]O0>d&0=ED#P+bXV=/(
)AK1K;_(;e\E<(\+R9&\DLPM@@OW-b?;2=_MdDNBX:,6F]AAIUY#5,O_HBdYN/AS
eOX<Y(,XWN1X45W@LT.FGJ\XP]O^>@?HCODKW9]/M1:fgYQMD48IdB5_F[/P&2,]
<+4HeO]6&Gf.\^16Bb5VD+J.,dWeDT^<bQ;,&gL)^Af7Y/9Af.IW0Xf990:57=J-
gX>L2:fD,cZ]_=STN=_:?7ba#A-GSHf5Q+c:UYT/41W8XWV)X7F9UW=Y?I0f6-Y]
4T)&&.6M5d3:3^H\=90@d.7T]YK)/H.a]7Mg5c1\OS)Y:2b63Q.^GMK+KOT_F<I<
YD5dB#6R,(FXG[Q-[Lg>PY4M],55;#=-VLGbD?NDGD4.fK=S-U5Hc--GVA+11a,R
_87gD5a?>G(N)A)BBJ.bR0;NIe\44Y?ODGV:W0W<BDCEc_R#OV+P/^AC<5MRY,&D
.df6A>_-;b9cF,UB#IPM1#gZ@aCR90b.G(B&N&=.,^aO3;C6XF1?X\=6&aYDIGA/
a6#7XBP-]HA-H99CU2fdFcd850PZ3U]OAI8O:-=(1\<)3]b+DZ;811]4]O#Tc\9_
&81Q7gV[D&B6cC++5?#IXH6G5:dNcRI.::\Y_[=4VccZ<Z7(T:Za-2SXX+\<DBP&
X2CP<_1<b1WbCQUN95/H0ag9d3V,J,/]DCg>4ba0@<S)+(e#E^/12-.@IP>b3[A0
TTCUSW_bJ1dF[U]AYM.9aMKaEWUW7Q=XBCLBC5?IE9+;ZH_WNbP>BGe#S+UU26=U
F.f94g2gH4^Qd9LBD/57c?Mbb#^a0cPYD\7^._VZ],,C-<^E-b8LEBDC_\gcNd_W
-Q?N-23(>ZZNEeXQ=4GUZJ5dP7<YYSLVFOVC980#cE-b;6WPC:__RL2Fd+1g_\8I
<@d\H06S7e=F(f6fd5,0=;C_M<DLIMA[>ZY7;CCG(\Q]BgL4AgFQ)RS[dOKF-ODF
<_b/c2-)YJZC9S:;O[]+IKF([Y0Z\f#^+J=c;:RG1_\NX4T-ZVH^EA2MQL2RY4]G
DYf9FK1K=gSab^(ga9GKa3:P0Z9HP(5C,I--b>NJXf2XBELA3_6Q](6d9UL:P5;(
VT.@2+O1f2Q7;FH.MZ#V]M.WN_OQM\1P00>M]2XO];QX;[8P+P>9\(QV\_34+SSb
>S+UX&7f#Pa4#J4[9/2FM9TGQ-[9/b<#:f/Ff_E=>=c,7Ke?>[GXUYR;B7]TB>W9
7&Z[08fe2gJ1SaFC+G25B1+#]X=BVfa#7AB:9;41#&474)I=E,d<(H#a;[]S9,5b
37T@=Dc3\EG>Z_HP52C9CU1MT1#PS3e#/])GV^L4J0QJLZ+I<.gHd4)X.6Vfc#R:
^B5;5L_/<4fP8cJEHM&D;#Z=Lf5M)XH7#4H@b_(^<@.RZNQUFgRTI,N6)D;9OK94
FBY6AX]DMa<G[C9^Y[I?W?<gd>-2?;cX9#CVZBIB.S^)@(0B6J]RN@TAR7V0NN3Y
a(V>d?>D=MW\C7/?e/-Y7::eRGfQ_[IUG6Ld9>-6g4\TS6IU<_/6ND4V:>9a>?<a
Yde4A#cZ4(Z2>1B#GQ;?[,Me<:,J#HbOULTCb6=<bW;G=.3.e,/3+[g6\IF#>V,#
(1Q0)R4_>17&R+POJ4QRT;1,Y[MP7I9-c621Z5Z3IQSG,:f&II6AMUU1bKfI0325
c13PG@c\JJ@N1(.O=)3A/)6ga#&g;cN0I38=/?@UUA#D7b,SS:-AIY@(ae(A:\>I
Y8OVTKA4fVP9,>8JEJ,+&W\W^Va\S.=#_7MR0-Lc(<EM_GW<K)^[G[2]BT_._4AP
X9WJBPYMB.I4R#N/]^6-N#Z^HV8AH?6=7.?8UUH<T<PI2\FJfZW8NJ/>JI@5IH/O
X#]2Ed#IRe[TQX?)YTDJ9W4:FX9GgW2U;P5,97K9[FS]eCSeS5LHQBU].]_@XURH
X.6OB174AJe:8bM#9YP=BKFI-J])4AE:NOefO(GB1DAeB6TI3e;B+:321G&b9IWF
_0a?JA+?/(RQ.c>O@(C:=;.-a=8(2\M(+Je>g]P/GNdR;f:[eL3R;#b0DDa5,Y)+
@N,eU#6=R]J:8S0eaU:M9PG]1F6[F6.D-#(2<](?\VPVI-NCM7(dC&#:KT,:UK.J
(E]NQ]SSBST&^CN>4GP,0gCY+2^NM]PWF2#E[A13gKX,:0548;FgfR<0XRY5#JGS
Zeg22^Z(SB(AYKU[(@2aVDZ[DW,X4g+BC1e6LEL9VS)=XaLIc#QR?59ab<Q/W&SC
O2>FYN&6TDEK[P/:RLf>JW^UI?g+JZebR^A72?&E^dELCJ@\0_d2).EY3#^bCCCA
5#(F3P,_\CV:X7Mg,5WI.59Je8W6XMZ3YTMB1K3TSU/5Q&BABM,L9_Y>eged3O)G
G8e@82QK^HZWXfO.,X^NE;KC,TgTVUW5=83EcYT:C/,:b3:34^O?0VeB,GHPcX6O
+L0A1?WE6=FNY=A\N9,A3=Y[LFX4F=6NUbL@c7_7Z4d;RY4a8Md>0KA>c_?+]TIe
e/e.;>\[_AW9:eL@^:L&W;FMR8Y>O?>Q0Q/9S3)UW5WLEeQSLAaD05&b.>KY-]C<
2FCZJ7T@]C>.S3bf993Z>TR3S[eZX39:E;[[N\A?\>0@_KPL#GYfW8UHTPS#M,5-
Z\dHeb4cc:Y\L+dU_ZgB1^N=K-_,ZR6#21-FUba(TfMG+)G=DdFXU1]MIAHJ7UU6
7,[C6N^2\_:7N54UfU<+APEd(Q3JZcR<@>G4;G,\d^V\^EEQ#3dK6KdR_#A<U]Qb
73)c8.g9+-&+dDe[>D1H-R##F>@[2U(3Y,g[P>-I<1DccZa8+W.\6HV->\X+SS4T
H7;#L2^=5WUX&U80^f&7YIM28=Y7?VT?<1(EN2&W5X?N&6G?ZLV^29P9E:IWJePM
<Vbb1d;^=0@F0(N5P>ODMf=^AfD0R01CN)&Y_W/_+gf&A5bY&,_e3:C;&;5//O@0
S0A,5SRf/b+R)X)<PGOEMBE2>76]e^V8-]E>-8M+[&B<,4]D:@gE(EPBZe;/_c#c
RdJ6aeY=GBWE4K]<1#ac\EQ@)CO>)&G:\,[]#IX0(NAWBT(,VOfSJD];)X)3+fCB
9g_&+QX8;.@fFPAR02L#7EDEeCOIGdO&=JI?gRF>(]DPd6?\,8=Y@]PC?^6P.4@@
6CJSM@O0/T^23WE6G[GO)4=GO0RJ.8OR+]JC:]ZXEKC@#1K/CegbNdc0UEEL=-&)
-#QLR/.N0gS;1U1@=\&Ud8S^#[L9HP.@09HfA\TBZ,aJ[.[V+=@YZG(aYBEN)I.4
5L_W98[U&&;A/Z&&O\OFV#N_YVf;/M#ZWgT1R,Y(PT]FWLLSY&ee,]YgSd[+_MP\
-?<SYb9;^_&7\7f&SGB=?(\c5M0N[&+>SZ:0CJbE@fA<>S.IP[FQBMZ[gO>1Ng-W
G/V&&2Pef=E:SaU4I\OQ>OOUdY8[(R^&LM7[:=;J,T_60cBGD:b\BEGQ-FL]Wf[@
f4814CMKJe^^Fd\Q1>BR[d@E,Q_&0,&0_&T<QP.&O@J_=AAUC8Q@2D0Z0L2LUEHB
3I@/S43Y[=VZ)>]GYf7fe0>F3f^e&f6QPIHf<(Y\IV@#]T:.7EW7C<IT\gX4-U/5
aI5,>f6cXD(KbeRa7<8<C4cG7OfRMF;LHcD-Q.+1SdI0J8W>C60dF7cFJV.:?Y>E
b5HgWX3Ic3Q>CeF<=+H/<-V/8Bf]T<TY&49g.5G-V9N;SPR]dRaZLX+S63P>@P:#
BV?5dJ8Kf>L=U;AS<;2YCY7I<ga\-&6J_cBf,PP<OK6X1=gS[Q9^(P+/876DKHa,
>>,-NE>9K\_G])18],_1cH_<_;09K]D)VOYSPWRN]8>NP#L3OU.L3IKBGXfJ+:JN
e>]7C<N@OJ-&EPegB@4C,B(A5C<ED@KW6HV]RWG(2d,c3I]@,Ab0(<I:\@F6;UJ]
##&1<bA\8YL5a[,D5bL=Ng&RP^;1;.)BIOH;C2Fd_NDU(;d]&gVQ>?YND4>J=E1X
-c<d4EWb@<X>@0TJ<2AC(JR+e0>-R.3B3OVV8I6J.8<1N[?^8FT5I(UATW9AG8#0
;SaR/JUScU/^1=9(>aX^V2TU/T9)ZQD70YK74e4/6X8)J[7REDCSK-b@@Z_ZHW(E
A?fKU@#BY\dWYS+0MPP8LP(EUR<<VC)C:H+31;>=L[e_KOF_?a<9b>6^0/]Y/1(K
AP6REa0P9CQ?.e-;_X?3AN?,faEVB^,,_,J+H;b(\H01P:HJb?:9AZQOO:6>&)d7
@0/b=OPT3/cOf>HO4WeOG]@9R(N^05,c0]B+SI::=Y._e+35OZ,(1b\U7K?LCM,&
9fJd>/Ic5BAT:34(K#X)Ha<@XfRMf(f:B\caGGUNO\9ZQ&FI&L]7aH7RTBNY&#dB
JcHd>?J1B.-ba-GDdP&O;S-W,YFL_G[<Ab99=G#C(4=W&XQCg<G?a?d#;<H/WMc2
X6L(2B6KZO=4I0<.78C<K&GZ0>-T(Dc&EUd<?PU:5U+A1=CH<J>(\.Y<8e(]QcLE
+\O)0D_(^BOES)BGaAX8Q^0R4J.@Ef;R^OW2;-18:#_R;ZG#3AFVYZg<LUgeF?5/
=e_4HcEdUI(e:9497eO^1&1_H##(X<65_./e2:f+;)^N&>7WP,-EOZAcFQ8_A&8T
a8)IU.C.>V6),HRR3,d.IJ_FbD);QDLC4^1^@E9Mf0HY1A^0aH6D7OKH>GfgXY=S
W;FPZ?KF^bFPD>S:9XY)/@fF-E(9AYITQ(1DGQX^71(;R25A-NB+=]4EQC6L_2XC
PgWV5#IgDL0OFbP0PFcF0=Y-+fSf-KX4=VN]_#.095F//DN<@g<?O=;ebPd8E?;\
FfC:QCT4D1047F1J8M1XDM;38;^NISD0P&YK@:JLKV=+B=I<Y.d,&Wa+FT(fI34<
1:[RI]Y1^aSL7Ef;M&.b6]>7Q5e4M+GT2U:(e8P1G22O:XP;3KU]O^Xa(;RR;/_2
ecCC(df&aL?36+Ue,TGJ3R@JQ0AK&/-ba:.\d-_+>d#P[7Lb]XV=eT_.0>a7[cg=
-_J?adf_KK(P?gIJ]g9[J4D?=(0=b8&3Z7L\;aOTV0>;D+fK8J7cL>_bB9XB9=)?
Oc//;3C?H<IAM;4+;dSK;1AQLQ+-15ZQC66TcV4<#4PbZ0-e?V/59>&:)C:FJ-71
B:JQ__Q1AZ:7RRCXN@O^A=<&eI,RL25T(R,3RWc^e4=7O2C,=<#.6ZbIZ12XAI,8
G=36DKP+0TT]Y7G-C#g-UN:)8LQ8&SYN]#>SaW3F1UWN#<E4HdOgN2U_[1-H=CXS
g[/Ob8.<B]42T4,(^-f.VIFNfc2.f5>GW/O9)8+<=M:[T7^2.MKGc@^>TC4Ua5La
/b^D)GT]_U:J]K\X1A)>8MCfV01XZ>NOTM.ZUe#MI1FN-:J,d:F.aa?0OD<T(G&?
I.D-dW8IX7#T@<dK)I8;].?42Ogg+P&]/EK?BE^5HSCZA_K^3>acRKdV-TL]a60a
T<1@]RS;D<>9&9@5+ARU2gLT9gZ3TI-:>e)B6X@CEF?EW1?<IT(44fEc3ZZK;g>K
d2CUe8@3Z<_#:-.9I[IKI[7UD=6WNU7_#4D1,b.6GTa<Jc2:@++e&0N?YYDfVCTW
@Q+@9XBRD14FRRW1CRKF+&ZO,<(EUB;_Q:WfecMeceXGOGV4;]=AMSV?g^3,4e>d
^a:_eH1^:-]c;]K[7.A<gUaTJ702#RBOB7MSJN8^\IdO==/+18K,a8d9BW]gKAKK
Va&aa/T8EL)W?V;SUX.GP@VXOa3VC/S+4&JUfgQB;;G#,1/CSI?0gNRB5KCWYC6P
#I>??ZF0KKE2NUa/(,.f4aI2L>Z=VZW#Y<:-_bF^781T)e##59d(?ASV4K>B[/+D
d./g<ZA=))gT06X^-PY\0g:&?\#M2\=d.75E]1683)+7bK/\6@/:<[U_><\Sd?gP
+<<eR(NO)F/<1@]GS@DUY8FZ>&1K]N5KD9[aL0LY\VK/?e@KVJPP)a5.PcTGA?,Z
,,)=6H#1.1J5Y6+@@0<<(X>bV/e_>We&?bKK)7B7g(X0Rb(\[:PF75SKg]Jcc)MY
PYGg&)L&+LOZ+AS(c:-d+P>Y1T2+2;]WDN#6cZfBLC6VgL=c[@Me#f)(f9:+9C3W
3Y]=HR:D<Tdc93P4M=Z0(bH59eP]GAK;70BO1e4(-D;DNODd+=MQf</6>KObf8/F
N3YQVQOOR[ePK>[)>EG4D0.4S9IHdAKH&(gO+e<<B+8NTDa5])fa=UeRaG7dF[-.
FPXa+g6;&VK[=]Vc/T7K)WKJG#CTA4TT/,(a7HJV]-Y0)EZTNV2NMI7;PP_DBIYD
A+/<QZ5+Ud/]-K^KRO4P6dc);KVK^,(^0efgM(Z4_-6OZe1gQAa=Q+f]d9U@Qc^S
C4aJOZ5_&A^CHU,TDHWTb0BaW/F^#.+<\V/N^>1TVFS.:/09>?&D+ddAS^PC7PDA
d&FHb:L<1YfgQP8C)VR@(LefW.=Z&^ac#,e:Ddb2G^g9X8SY0>g7O>T^XY@IcL2J
JKeaT62MM1_>MHV3\C&)>L1ZRW;YcDY&Z,YZSeBN\?G_\KTCH7/3Ea@@+BMI&+[a
F;,)g[\6R5X7[COWPAHe@JS3(?;N,26(?[Q;BWH?f-\=&gg9#T^.@d+:K2)/PZ)Y
+T=-aJK.EOE4K9FKeL5.Z#7OO:[/M@VK-6e?FIC+c&[U;&05eJfcWKXJ2V>_<(V]
S4JfY([Va6I#>fc+HPf/WRReA?I_&0W<GffdPA5VM#B-_YSR3#^4S>8W=CW-fWde
TKGHZcW&1XKBP6b<H[;9+YE7-Nf>O\NKFP@O\9=gBFP-YBf(GV]_AfRM88.8J<58
NW?^G1TNHJEEe;/+)GR/#1=I;S8f<T?+dUgSV)_M:)ZJXCF:fSGd8eZeC2(Ma]6[
64VR1DW+V,?EMT>VaLU1Q/7WCg13H[&AS^d;_&>0/c7642g03&0O^/DV:8O@;,E;
U:aS36F:6L?@^9SKLaC,S)DVdWZ3dDDc5^Z=Ea8S;,P]ABA68RT:BT(]0+I[0-c6
M_QgXNT86g]SfgW&c8GNT.U<MFN\&-+:CeK:;Mg#R0M+9^+=^Lg1eQA-HEc@Qf6:
U5gb4RV[b_D)XS]A/N+)+aZ3O+8,-JY)bg3]2=b:U8XYA^W7JITF0<eD]BWfa:DC
R65?=:#+-/3C(#R#/5d-C;,P<0AQ/Wg>SI@)VN_L(S<#_(4U=26&IF]JGOM@B(;0
fT+fRF-C8;+1]d])1;Q#bF^W,N0=]WE5T]82S(2@b(?SUcX=Y:[R(_+5OLc&Mf&]
3a?@3_gXgOIYJSK1&C)XH]FT+b(@-MI#NQNS<a=B@19^?XT@Z:5WMd87JS6^N>dc
ZT+5>LEU)cMSCEG_AC9VaNKDF&H6#H8ad\]\5M:9YOYJ,5(4ZDL>H<eZ,@b:J-J0
)?EUXI<-;<VdbBUY1Ob?,.C@ZP<KZH5:3_C(.\GR;@(R.K[-0FDVR5b^R/FY+2P:
91Z[WG7]EBJ#;6cG96N]+;NN;7/Z;-LIK<6:?F0NgA<dO4U-NGAa.T<)3P/_FSN\
G#CECL;.F[M(RB=U0Q&8gJWVBPPbc:WG,?8I_<6WB)aOIfb^C,6AXEc..:5VN+(Y
@-V4N0d(Ef]EQ#7a\7a7&+Z#Zf:P#3&XbL235e+g;O/a8cRE?,?,6&].4Kc-a0>[
ODHF2Z10(4]dg@-gfObA0,6-4=C/IF_L>&1;XbKOfS28ZKT\72(X2EQ9/_+a7aEQ
dE:9#JUG,)SW1N>9eO;)DDZI)35+Y9.;^IGH+1-^f7f+,57b=J9E2N8#:Se(X\A,
,2#0D2+VA&.B]0A@?g[-1P9PN?DKa1GK:K6Dg\O0?Q6^BaIJ_R;GaPg@WM5AccPT
?Fc^<@g:&cEBLQ<\GB4]2g^b&9+a#?(TB9)AH1/=FZ1<Cd,CZ(\FNdP@:e,TC@)[
]0;O;e)&&Sd<5Bd7Q#D6G,dER]KJ,,cVZ<UcY>]P;gc)[,]?T(#C&GfJ4O/TFdIG
&L5A\K_LdJOE?Y\3)7?O0AJc=2NMf]=U_Wa\<d4c(Be,UTTU5c[MZ2;2JQH3@g(<
MC@;4TbJIV()aeU^ZAYQ#aNXRc5ADO.ZR<?\FFE(AQRWQOe0(Ha=IP?eB;2AAd=9
YD,J6-b/cM3RCK#SS^U1W3J2c/J69_;14Z+N:F5GgN?B>]Y<McEWJBe-R)+7Ba95
bAPC.2.)66VNfU^=)9-0@[IHIH&[]D[3JB9PK07GV=TD(N2QXK^Ae8Y97T5,9BVR
@.8U.6R\WB/DeDPNU1YS).\1I>Z,HT\D#J6Y-,0PKYLac_5[+FHSJF<.=aFU#:b=
SCVO>PO>M+f,de:J@?5@K?)3d6O(3]3,EMSR:S@-=7G(_a\c(7F>A0A::+66-g8D
9JG8+\,D(CaSVe@;=0(f).=18]&39<K9P3O5a]-Z^9(A4V@a&5.;OIUV<UJdP6QV
WP\)3MKDb,Z;eD,KBC6]R6b0WG#_NOR\@F?BB=Rg&Y-KE3C^P0S1I/\P6Y#Q9?#R
/5.W6T3Od=Y]d7eC)U0E.Zcg^]5</HN99f\^bQ&LOD<3FM:Z_8DBI=)JW:GW^U=+
V,fE]Z\fNfMG?30N-<cM)(9V)E(\K6F93U?98ceN>60IUMd]/W\]AXQ+@92.LJX)
DRTa/d&0ggMg:0Z-5?;3]E(gR/X0[72\N#YY+_&aR>&?#CFM?=?@-Oa9dScRaP,I
#8T@c4GP8a1P?^4+?X6/e@>(T&LWCAfQPe@F[.R(CdN@37E]BB?^VQMfJ;C;D1;@
M\Q27Z)^E,#Q>L\Yf,SdK/g<)SGgTRHbQe^HWZC0963FT^cN>&+R-[V6B>9OQ@[,
TY1B;^#18QFIg8,D&N=LZYV^@^VV],(fUKBgTL<=BgDICOGf1cANeA-THA7GgK;A
(8@OVE5]2_-SN)QDO<g-OKI^Z8\1K[d)V(I(f5>CJ@YOg5QI;&U;S^]&4a[0?N8d
=]\b+@NBN#_\1IOeV#ASXE3@:49TJeL]\)YZ+F(2:()_FZMP#6#GaK;@M:@V=(2Q
-=VZE_\HEgTI8Lc^=98,c+V)13T>G,_G6M8HC0O(U6B&5a3@2T1=fg_E7=I4^2]#
@=FXY6YNA_Y,7)AF7KVA;g_8+Z:D:;,W>Y6#da4VdY(IM&#P49H:WM3Jd1X_WLV;
6VSJVe>6BGEMf=//We&AJD^gN\M5a^LcfMYT>P96(1.8=TY/I.UU2FJXROM03<H[
MXG[QN&]1<eDO=-@IKJ#fZ&-aQR]AI9M6@2YgR5HILL88T25=A99E=W5_=Y>PS<6
c#[K[4>7e[S(APRPG[P]ZS&H\[3ZQ^U9TY/^0df:5W<\_Y>M46[0(,S[,Eg_LXOH
2;R[;^2M7^PaK@8Z<7<SBLK+L3/dLRBP0I_56f\0J0@3++HKTbgGIA&@/6RFVbgB
P^SV#bVV#dJ];ZVBSRTb,\=\WPW(;Y<(5,IB(P>PV:=L59<)c;\>GD20g7U)U3P_
g<3P3Ca\9Q/,5d-NJJX+M@5R<(O;R.2W6QU;GZ#fP(;^<\VOg;KZR4eZA7=JKCg7
RMZAB@W1)+-X7Fc7a:RJRE(f3X?@b,2#O2^WLg.=EM#TB_09[DJ/\(BV:=C&cAK4
G92^(G8-W\>B&Z_TQCN;LG[MI#dIJW&b^ag2PQK9]de\8:Rb[0I,6U;TQ4-UB#,E
7_=UPX+^8VHCc/5/A9CUH0HMPF>Wb8@DM38R5Z42\8^Abe304XgdRM&(ZIe72Bb,
3#[8I_e3Hgf#^S)e7T9#0f][K?)NfBKB-=))OHD>2TA^VA5S=0SH(Ob^SdePM0Lb
#>I=TDKM=2a42-RdX<QHc/U5OXfQV3NTf=Y85MI?V?>JgG09LX)L,@G_C#D>RR8U
NI.OeMMW_+-PQ]KRQ_B7b@\cL-EOCU&&[ZQLe@+<6R<_9fA:?-WD@UeAC@Je(?[#
<4#E)g[1-H-#cA6@/Qa:K:ReAJQP;)TP_O=PDYP32CVW0bKDR(_EAEg#2\:_WKHH
GaXDHI^^J77DRS9;\K@3KMA;PBKYKaE;BCYQ[R?#XY.:.ZcKNF0Ye4F,Q3)KS5K^
IAK[fQDM>QO-A(>V<P<&6E1IJ9fRBeGZeb<eG<3ECUR;@OM?^@g.)]^O1ASXJXC1
Z^U9bDL9FAXJY,_>2J;FFZ.3:DJb+:g&_WMA.E=U.6a+E9If/)d)0+Z<U4TQ67U1
A.?Q\T-Tb+&J+7Q6U(Qff#78g(B4Z;NO\R=H6:CL8(E,eT[,WXVc2U=)7<:cbVRc
74bUd=Qa>f(E)T>MMfE?^:Q7YY+GRLQ&M:1<)Z?X.(N6OZRF=Y^FEM7,M[51-f^]
e6TVVF#.J6J[UdI0U6gCE/BD@1Q#gIUMab:J[L3(g/&#([,dd\+(?@N><<_3W)?B
F:7;W]60CS18EI_F1fa]].Be=f@bBA)2)L_&YeUfI<^EE4ZId+?aTZ8a>O6.YR=]
(5&1fDW))/:,?Q9d3>>/JZ8K8e);5:Z5+Ra+\Y[Ud;a9Z]N.IX@/c+)=Ua0eW]W6
]YgfF&#+0:GL-RG>>BR/FHFCaQCVe-)68=3OCGV[)V._0[^^GSL_#Zce&+,)2V?L
5^4LZ=4IX:1Z0:;ERI[88O-Pb,]#.XL()YD43C\9=/ZS4U5/aBd2))4OZ]^^1_>(
+B.ePa;FK]T7P5_ee005f4gH61=fBI,Fc2,\[1N6S@(:0VdLZP^^a>X^3_G[U+[d
dUXbG4QCdOGP7S9Y+\N8-^8LT,LP^Q-OFX9?9TW?8WJ/SDgWQHe;Cf,?1.#+^d7\
#XJCPUB(1B//:R-/,=MRdU,VSZ&&8dJc7)9D^cPd+geYIR4a)a[TK9b:HC\HaKTY
U^f&_CR]5_<P,abDILSb]/X(Q:RLBCfX#_Q67&C]_6<#g,f,.EFO8MY#W2P5U8FT
4:AZH1W1MDV>N@JRUd1Fa?=cG?)G/-[@(bWSVe2Q6@4?DR#V7f]@E.^HUJ8CRR:[
Ocb[37CdO3acJOI==Q23E,M;I?1U)gJT<c.^eP>Nb</f^V#c^D#LWc=BYJLL4@#b
VTBPA:OM&DbgGA0f16&b^Q^NQ3OH;J>]EbfZ5GT,SYKYD;:KfR,HUDZ;\F2ZMG38
a2(J&.=Zc3K<&=I4_-?=@1</A\YX95JSP8A7Z95JGbS^Q\Z.?M6A@Tba(<.e0RB>
F2P5DE8,g-3aKHeb[bO3@,P7cLOW,@E#=<5^TA:FDPY>R.<SfLI2c25\)eN^3b[B
BPUc678Q+399M3K^\<>6^JL,V2=2Z8cE.MRP?QR57Lc9JW)R\ZG&Y:3:;eWYM)1N
]1TQD6@-^J7/5H.JT;=\C-b^c0/aeIdG#6-EM9;C?W6>7Q]OHbHH#Bg2=]DS,?Q>
,(UM7=e=b,6V.K\&M?+,Fe_&AC+CCF(RYgGIfV\&LD^\+]ZJ_L/C)E[@/4F_;,HP
gO>?)(\Rd?QRQ@0H;G2a9_G4;W6J0QMQVTa\GS+>O-eVN?=.^RYYD7M>LN5O:@PE
EWCX&=4GL)IX^L>_[^S7:<A,13BfUZ-.6-I]PND#TgE2ae+H4-SZ4<U<X^ETYBc.
?EI.Q]U;=G0SB7;36J\4.FA8Z\G=&b[FDcAW;S8LBcM/91K0MW?&2e\010NP(]eV
@7148[9N-T2VcES/@?KN,53A?+M7894?[,7d2GJNXfTbd@G1TKS>fKU4?WJ04HA3
4@7:Z>3e)(W9KS2R974YEa-GgNM,19T)AgOSWWJ>&RgQL_&;d:0D:FM(T&O.M9ZS
_C_U2+d)M^1TW]U.Gc>TXPHeQ4VZNf9F<N7/843EQW83:C03aY&T9Mg-)Y#XPN_2
N/6I@B/9a56Ja>1\U,eH5L)UQG3]7MR04O/NJM,1b+A-c@U\MVJ5-<0NcKfK90e>
H<(]I^J>+>SG6+-P@9\bDeT@J,D?>LI^[bG77>9E:/<eA0Z5aGC6<35#W5:\dBQO
ART=^2M(cA3WdSP>cHY(C;<gM\UdLeaFA:Ia1S0J;>/Og3MWG-NL?[-(^7=LdI0=
4=N=WDa.Q/dPO?)JC=U);;AT:<9R&I36/CJ+>e2/)F>0>3+38R_0_ec_a9U+QKVA
cM9^:YdKEE[I,Y-RGA3aX=F]>(U.Lf+c7aUT9#FA,B<UQeM0g<:GY1<U7QZDId1U
[,W)8T#<P\ecJ.6D9?bLQ1F9&HGI<cD)c9UU-BI#a+L_d-L4PQWb;L,@=eSFO6L\
63X?<J,1ZJO<^5B/e@=84cT,3dA)6>5T1;Y&^,1#Z7.4?\2ZI;P(#Y:f20NMD&?&
QA17Qc9?:I]HEUGI:O>.XNI6BP^+AYU+eDOccD?-+(D#e(=B.0,157YYf.g[V]OP
0BNSC:[]W)@eb3/)IL?IKHcMILUX;OVA+ZLIV:(4F(d/>QFR&TQ=;:F^V1c:DV1Z
;>gTM_&:MC,Q6B4SBVQ=5:a?LPTU--T=4Q+HVAN<E#<Y:G[Y4+:/C<#[O-Zc&#;9
Z^OEE4[bcWDJ3.MCQ1KeAOQ@PT^D/6f@U:aOdBPDJga45_#/HMST0]=GQ5d<3)NI
ZG1a?5#A&9D]9C+<_0[26YV_UMVHf),+f8S)X_&2EId,9TWC8,7I#Q&&9+,1]IQB
RS>]NY;b^908AFEb6;9K;Z;.eMJ<f,V[ZTJE.PWK8/@AbO;H13JS69;MDAN13@R+
VA?6=c&+IPUI^Z[<?=>83#-)2BJ<aNFY7_f2V38^]Pg0A=R:ZGCFaCD9Y>aHSW:1
;[@4RYRcD.(YAUCF6?PP/+9J^Y<QA<QL0\6?e][Y;)YEL+#I4?S^6:?2W>)S\4GQ
U8LMJZ&+T;ZIOX>EWUR0E&5QNgUYQ#SH?@:d31A:g:[;H9GX>=83[_7[@Y4FH<:S
XDR:HVIb:J1P5.J^gacLcD,T;&E&,Ld6],;8XHJf;e_a,+&KE?9W0HSFRX/>a(I#
^<50P=8/=c5IRTNIb5N,1O79f(.BeO5?eO)^D7U.:^>Ta?JcBP]WQ#A]6ZTA(gFY
5V/=DD&(&YMA64/S0I^E#Vf>EMBYZ,WcBd-10E-[7<CUMP,(Q2E/b]T\R9ADe7KY
X3XFIL6SG8O-^b[U_eLa7H74A.R83bUQNK79^(2U.N1&J]3(#I^IAF=-d)+QCNI^
G>>G@[#K>)]Z;>2ef[M<[E>X5Dg?gZNBBP(9Zf#[4743/>Q8^ZbMgaAFC7UV:-O8
0#(6G9NO1W>5g4bIZ9(COc+=\cd?/+V]O2AeL8NFHeQOBC5[KJbZ-7Y+-HOW[X)D
fJLC1SS?4Qg<H6=W;XG>6Eb:(ZdQ<^I=+-A+&+5(<Ye<gO&-]60^P.+:4>C@W36[
G=-:1H[@#BXT9R(AeVbS:6Ngea^P:MZ?D2eaQJMW:TF1R#U+WT(Df1W_d3NT6D3)
G,<==PLF2KAgSLQa<Y99=:VMFaU3E^f0&4.U],U0@BOB/e(RJg<MfA6BG)#cOIOQ
#9H^]\PJ:DM731B\-[HZF7Ib<ZV0N>FAZ=f/;9TIVRPODA^?O#VC(;@,Qb:(297Y
=6JDYa1\(;d.4#\C?.F>(2,3D\F,X5K[5RcJAa:NY/8?H9f&@VA2@VSN,1\f3d^3
>7Y8]FFM6DP;;;CPaa9,#33[(N29>)<.BEg)UG99W1e)8KbC:]9P.8BcT8#@DB+N
K#ATK/--6FKSgHdKS.Z].O=[1W>SJ[/J@dG)10ON,Na:e6:8IQ@2M)E-fWB./-D)
NT0Bc37UT&E]R@NdK9/^B@NaH?dDQE[1Q+M+@42CNJQ#ZS_9YF&[;\dK&&P4a[(e
JX]6ZNF>MGI?(f(A4:)EU5QSD-aOVa>:6>4efB_)-B([_91C.M5bO\1<<#-[fY/+
EDWgc=JQQ41KLE2&H&0JT_4I]>1OVHeJ)O-)(@J4g4Z]QDYK\A5#a>7OHK_#&FaE
KaBOOBQ=\FOg5e//KR^@_PD1RI@2I2d:e&;PM<H/;Ggc<,T5&+gSV3+:PI^BEBJ^
FZKU6OK1W^?Ef0Eg]-4VIT+5.#d^ME.fVQ9GNeI\)?>H3UTFUN276g/4/Me1@ORT
-B3?6]CLb>W?NWLHMD/7=_(O&O\_<>G#WP>IV37]C,ZeSY1W=c?F.N<,/#4R)aXS
-3D]EG)dgC@gLP&Ub+cUW,aOS9/gaQe?aXQA_8f/C.=/GFd0BVYRb.^DAYI1Xg-3
JH\BU55Y#[3-c=CZO8@JJe[\BIN03\U_]U+FWF)W5WMBf5BE/B0V#0EC(+2\:Q40
]VM27g>ZI#1;]_e&Gg<,WAE>8Y6@4A;OV>a,XBSca88_BU^E?OXH-SJ>bH)bOI/.
A>/HC38GMPP.J/KPf)=eC9?Z=O@R&^GA)(]J,_LK=T,>dJ2^/[a916XHY6>N]&g;
gK_YcS#dP)5];eBHW38(MNgV7@PW4X/FKMg?HQa9e6_(U..S^1ASW;&g@BQ-WLC5
4<4(bQ@,VSS4JE.I:7P10D=[3>.d]&L#U)eOXFMWPQ_HURPD6g2:+:dcV-6Aa+\b
F.#2,&FOC]ACe4Y[^_<H=+_0SW#PUZ+Y7+]ZAW?:=4V6c7MY4P_dS?(fg7J(XW(+
G:LcV9(JEQRH.7beK\SFBbeeJYD>;4&J@g#YFB>UIO6U+N4cG5]HVM?4GPV+\f.e
V[2cLS9F\[V\gWB(DB6>ZJbRD/M3L#T-XIMH6TUW\07fa&;c8,I3]IKA\CVF?e0\
V4<^KV,;N\4IV_))H8(I[G9A4]15HBS31<g-;;^.KcKeBfW/5aLbaC5KYO1<\CP?
aaQFTCEgBeKe&#BC+,V>F\CX14;0)b02c.TQDI#8PCVPRXU3[UB?Y;+(eMf5#>NV
8-_S8=V4T&W3_b(@6e]P/<e;?eW.Zee[e8;c-d[N/>bH1XE&BSLLb/IAA_f>>78>
A3CB=<W#Ac4b@Y2/YJFL2->S8ZKbZ9)#&=ZC=0AAX_IOfTWU(_Y=4=O4#>JPW,O4
1NF6^cZND,9bE,\8WODTJ>Y#6D.8XBf5QV^Cd#>0:4_L3JE^=H]06f9XPR+ZV;4L
BQDGQ/W,/;a^7?]cYf:]:=0c:;W:IYO8P4WaF,BJSB,?1,:+QA@88DZ5WaOEOePL
9Gd,d6a)f:>Z7Od.HT8_@<Z_G32e\>d>7Z6(PSRH?A1H_fR(-]M2@;HXZ;OBb8>Q
+^RKTPRGT)_,8C#RJbaZ(@(T9W_W9T(T)1X<@)<9K8WBUAAW0[+F#aEc7d9\92=D
P1G=81K80R2@5V&&BM)53E]&\E+d7=EP-C2?d,D>M^AgMb0-3\#g0Xb\FXMTBY:@
dS4(H\>?9/C:e2DZ>(P2W-R)]IOc3]Z0Ve,N-DbX\XPU&e,b(S/30a6O+\e^7cDK
HdgQC7QJGU@ZL0Z^L4EQSEa^N7^O0E(71a=F1FA?H#f3?F[W,YM7fFF^,Egc5_)d
L^T1D^Y-Sf4]OGLVE^2eR68U_TOV\I]P([KK/7#]@T/019FGXggJ4T50@N\_#F#>
:<WE1?<IO8=B&Y:(@e5KVE-caX8\X7CK>5[Cfa=[ZAR6>ETJcdWRVQJ9WQ<PG6EH
PN)fSZ.^AQEC.B/,XAA(QD-7D,Y;219[CZfbg>;8>A.6ZNWY:^)AE,23Y;SL.gV8
>aCb7c4f8AXc+WT^J+<[+Pg/?E6b4X9^CT/@>6XWEabSL4fI5(D9Dc)KfL_,NC)B
JVYe6S6Mb;T\1]8/B1UK8e=7Q8G/6Bfe;B:ZI_@6W2;]N\UG>J>_-2P<?:C,F?+<
U]Pg(5^T9,AK8D)g\.add9(-VB.gE][98(\e&b&Ie0#88)c5S)@7,U&T7K/6Nf]P
A470B?8:V6Pf;<<I\aTE<5-<8<+dG<(F49?)_]#WFAXFc,A:F.G<g7P4Q^E>9U/W
=@0P+Z-<C<:G#X,R)+,W,(7._Mg@2S3(fU-e&:KFB\-YO#U[06-,:Q&6\@-VDRd#
#]4UF<2_EGGN8-KFWJWZ=gJAU/1MRES3[3DFC5,E:T3-)7QW<Q&U[A@1.P6W.LO2
2@5GXZ<JFMcZRA>HU[);W^@SY/geL:gWBQZ;@IdaeEU@>+YfQ\)L35<Ea1/Gc/:H
C/3TJ[87+0d#6.\TW=[&A7N2b\f6-[#dF_gM19:8X9X?c>>/8^2,d\(]+,Y7FAc4
KX6X^&+LH=,59_b1Geg+BJ;_)RS-g@+]VGc<g<^_(aAZ7@G1FdL]-_T:AdQ.2A64
g7@d9[e6Ke<3Jc/N2bGAgD9a_>S0]^#)CO5#,aQM\/A)&fO6LMfe_J22Y&=JW/JI
e?>-LaP:SL_Y[1GSbHSD4Q=FR0I4SJAQ2:6)3UVcE=Seg:aL1GgGF)DAFS3gV=LH
3,DNKP)gOV3UEPQVbRFP6cD[g63.IU4>?IL7IZ-NL=&5WK;EgMZQMd^fT_.K[g+Q
+_eLc](Wd.^(CbR4002EBTLH54E1V0YKHdMa)f2XGXI=P9A=6K30O61XDEMBI/B=
NSMK0C(#\M&BG2<#JO2K>D7NIX(<CAD,&.K)4SC0[X,<7LWZcXcdP)6b-]J5E(SP
79O(+d\DdG/3]9N\,gF6+Z6\QbL=)Q\G0XKKB&K82Gc6[GZ&L^Ne_ca,e:V6K^FD
)5N<?ZSCeNKVELLfV[GX7?+bCHOaffI,P7V2<>R\E_Ld\KM/9ZL.[[(Bb+\J&bA?
T?GTIc4Y+/08;#^[9aVb5NU9A(,_AFVCZ14.VM17JXF&<OA)B(YaM&4SOD>:CRDY
=F.XUS@Y(YTg)SR_:+eNbRG(8L?X#)>cJ4+.X2XL]/g[0e.?g6YX6gX9[C:.;,=E
?gDe\,6+0^GTHH;J.a1;bcV5\C@/B)S7#-VYe];YS]S25b^_J\V+J0H.N\&1UDE@
4eKT#_^++c^RC9[(D<J,C.[NZHf07D6DD[TCeP@WD4aUSX]STf<V?0JP:eBBZOP)
E+3U,.@@>C#?:JPKG<:#8M[TDV3/:12/;Z7+A^>]&a:XLOHW1F0/Lc\G=]TLgTX,
:;>\SFTA7B87=YcDAK2]Z7ZdYP#;Ad-7a4f.:@a,7BE#:W#:C<4S0<gbB.fJR7:)
4_aBFI\Ke5T]491OJN=1d?M9.,-0(_7&KHf]4PbT4EI=[L<A?dfG1;JQPK.NRgBJ
G2^1)ea&dL3L+cH:3[LH>J+cf6beJ^f8P,3K&0W\Q2N9cW834Fa1F3b29&9POa;F
W)f(VR34_:7J9N391^eS?W+D.0C4^ab^3Z6SZW^QSc/CE2HdI5H&\6M9U^[IF6e9
UBRCU.E7BOfH&PR1KWTb1YHdN8)?+Q0QgG9g5LF_^5M17M7<-N99d[<>KfgQN2ce
aL8c;6P[OZF9fDZ==d:YEdM2CK>c^^?-U8T-R@24KQ2gAbC</0-5HH()Pa8JV.U1
5[-<0?QNM0bFZ7@7/<[6#/Zd]aP;TTdPIefX2?J-)c+IfJO;T,1b&,EGC@d_#),b
QT1@CFAR(-[_dUW#C2>@X)-,#DPJT8BV#4_a5e.SedDGHSI-7=TKC/419OY]6/_g
<W-SbVQgG+M0][FM_?<Y.P.(=GW\,KcL1L/H9L8+P\DBSOG)L4\e?g8&L_K]-UN5
52G5;GVZ3W1<57/(bSLI>d,G.CB7gX96SW]BSd/Pa#&3TO+E/,>V@50dI#=J@4O-
>V)C509C&\#WF6e,TXQeTJ)f-O#^bAO?C:ID21.Y.=J:1V0ZUU,UDfM,2JdJ1Dee
79?Bc[:MN2TH)d</-Oa@;)I@W1M<e&\LHdGWe/N\eU(A7U(4CELbWECbPfB_F,R>
O\NT:DS2#6,/DK4M\&A]&@NKXTfD.8[\e8@O6D8O)<gVC8Q0?dLJ>gEQW8f@P14G
N2[AU3F(SV?;(=0ENZ,(QQJ6ZeL04bX5L-EVfMCA;D+N9U)J4gQ/-[V+4OJ=UZ:N
N:&JIK^A][H#R5?4?gVK?K;BR0[E9:g\M4F(3.gRF4Q,[2a7gWb9F.ZTVFZ;^DB+
U,cV5AI>-52,=R.0W61T^^FUQYVS8Bg,Q;fFe#8XZ#I;=W1W5eRO=:>.].eHST.U
/5N(?)?[TH5M.PRQfAT;A&6Y;Q40V.aQ.8MbgVC38^2GfEVZ6F+cJCU04Y(W:KdW
/U-P.1JNKG4EP/96HZL^PLTW(Y58_L/:U1_bU;T+3-J=+FWJ-81]?KB=H1Kc28?N
..CR2&DLT@+5-H>:<-8ITMHO35XKB.dWSeU])A#72J7L/M7?4BJ9RHF#RCYB&2L@
4gaGgUbVAY;I9BZeK/,T1I[1d9ba)6HW7Y8KE.A;gPXLA@6.e7I>SQ/0IbSfM=FF
AcdXI-?-)BZg,R_\IWQP:cg94f[M<f^<C[)FWIg.T5=LQ?d<R_TM=28A-5cB?77X
M]4H(1GgUbB+9)2GYW1Ga2cH]ZP=VeBd-,=bJ<Pc4ag8.N<BLXJ@R,HC7_H.296>
ZNZ?2V&K[L<dbKI\ZMG&?:\S5O.4+)9(6-^cO71N;.R@UQY9DaLNg1=/<57ef\=6
16Qe5(F-#Le<,O,LVQHR8O:TY\057&\.1HZ75W.B.W8HATLHR>?e4T0KMb<&HY=?
L?2>,f;.a_7+Z/MYHY&6X_?6X_WE0\<gAe2C\K.CS9.#MV9cA43+Yf#=&;QF,ZLb
U@R^EUCO_<RBKK.9OMb@TcHDLUVD5d5(S4U7(K^4af9CCc=W)[3G)N#=I$
`endprotected
