//############################################################################
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   ICLAB 2023 Fall
//   Lab04 Exercise		: Convolution Neural Network 
//   Author     		: Yu-Chi Lin (a6121461214.st12@nycu.edu.tw)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//
//   File Name   : CNN.v
//   Module Name : CNN
//   Release version : V1.0 (Release Date: 2024-10)
//
//++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
//############################################################################

`define CYCLE_TIME      29.8
`define SEED_NUMBER     28825252
`define PATTERN_NUMBER 1000

module PATTERN
`protected
T(T:0<9/FRMTbSXe7K/fN/D?^#N(S99bOD9cWL_;S[BLB.e(UZE85)4XFOW^\L^:
GYX9TNPZB4S&/>G-PA,<VI-(P;TaPVB\<Q)PK]4?+XU:eUT1\11<B.dF/R;X20X6
:0&FG9a93VeQ]U/8=O=WOKZgJ0Jf[eJW0T+LKgGd+Q-<@:2G8N7UMR6KGNC.C@JF
B.C_;f)/C4Hg;PM0[4;_-7IJX2LfI0XQ-^D(GPe#af/FT@_fcP7gP40IM(<4(&JL
&PTfPP?#;&KHH3_1#QG-H],#.:+)GbEg@gTd^-?e[7b:/CHgO<3<<0DQ,)WbH-PD
:Bc<F,A+C2U7M0G;WT/Q@Q_^]Q-_U7bPcMHF\;3(eaeU^]48b\W[g4DW1=74E/c7
[0X7C(X3NKLHVGQDK&FL68M+COFdB6acGE4g@bgQ-g&/;DR^bD)LCG2RO=_>#W<&
H^]bfcB&U2_[AOSVfFf<H[.;:@=.R0Wc#bKS/T.K9M0+A;1@+KI3I,Y)#-M,YV-/
@D4Tg2g5abXGLLZFB)\Z;9=)V8A-VUO+=PG/<5W_eWVcg7cbYJcD-ZWW=I-<egf]
&cR#\DHQ(C7-F9H5?[KY47&EF;?/RJK>A-YDR_EWGV\gC2=VMAaZPJUZ?d=Oe#gS
a&.1389:BNK+((g=F[:S]fCEWT_7ba#ggIV.b@a@OAORe#;+MW_=a.4.GAYb:9XT
9K:94PU)G8TB?++RNN#N_\Uee=O?_b58W5H17c\XN#XBYL1\(^c1HJ]#/=GUY1DI
Zf/Dd_-)P1AcdFEW(K=9S.)e^<RAL2XG7+Nf58)?E-BJER#bKM@T.:VIQ/:CB_e^
G-0^4eLJWAJ;+\ZMN:\AP?JXG_f@D+P;HR+YaZ]gHV((=I50;;OA4F0-Yg@LU7SF
LNd]6a7)OS)_DOc<bD\-?]\4J1S>T-9WZd9-]NaAOA8X_;_G6Y^/_Ud6fW?D()OA
GSI#ZZ;O:CfdV;80HL.]&AB?eJ^)=g=NT\R]\H2:1NN(b\WZ[K3?_O;7W(@f_1b<
^Xf:=#b-22eB8d?>1@5U[U;1KW<A-fKb&Z985RATa?(P?]4+AaOIGWCL]gA.7W)e
7.(1;KR-<3^@4/21=Z0Ge-VOc4P@KA,d\[S+ABSf;\d<aW\52bfN9TaAI9-ETR?_
N;2PX,[5_L=[D/F[K#QV3:&)G,/38\[;-2cCJ]LP<4F??^)70OPLTWW\#VL#>A8O
9<TSgd38POa8d,aB9JLH[-P1JRL2IF7bJ:Bb[49)CJLc2d]=N34L.DO(-gC#)RM9
QSK.LA>;aZ9@NgSA6_-70^N,+L.d4RUfLW1QNb_PR;fFGL4NRLf2S_]J98/W59B:
H>]AP_d7^)-9ZOV]g&a1@<43R5WfYGX)6\Wgac3T98+/Y-UYX;=d&BXDe&?#P^OI
R+0_)YRcbcH&0DQRS@a4O:dVH.G+5Va]-(a<Y]OV\b07P<bXGVI>PGa.gdB_8)EK
Y:5@K,^G9):J]EII&<f1bG5BC4Q?.T5E];MK7K0WGI8K73HdVf0CgX=+2RREYXgI
CTd[0\BQI(&gK:MQ(N[_C>d3@(][I;6B.X]CE@&UAZTR96d-d-K\]GP+O5Id1dWI
-)SJUJ9cQN-2X-#g+E9b3GM@=UZ\/XXBZ-X&9Xc<?b9ZX6]EZJ^.1(5DJO=cF6@/
@80=/TAE-O_5EBe0=FLM)HF6Q8.J8)Q4A81Q?:G^d8+f)[?[CgK\\Xga\a]g=ObH
6[7S,1].EVLCUU@_XLdD^@Nfb=+77I.663\7_(PO,--c=\LZ?@\C)&5,;cYbH#V[
]@I8LTI@Kd/_A/8]c5XGN9?HPd5_8\)7CgT0J^1V2+Da8\T4aD9S>#V=,_R73/<&
\@&2581-Bb9)6F;ceJH_[]^5NJ238D,.?K)?6U=0F0&[dE&2[<FJ]2B/-2(OEY>_
0I;X9S[0[MEJ+8<<,BP<dQVE+4V-?Pd]8.#<R,WHbLIE@d.=a./g#E^7XT9WA4BP
,;#gJFJc0e_&Q)/,;7HcAL[<CSR=_7_EdNV-KH2QfAO]?9@5O<KI<Y\=8#-WS8Vg
R.bVTCfWX<4G6fc5AB,;g_b7N^F:C7;PE09-FI[DILZO:\.?6B@FG>9</QW4[+]V
UO9d+1.W[HCIWB.+C8<,S3H(5UH4e>eFPT4/\B6ZHVU=K/,cZ;&>V./3XLP@e9c5
[ARSd3_<\NSf5+cOcPJ>SS]#BFJ(75WW=MSc@8[J5]#[0-=K-]M.:DD.(AESKf+Z
,<>19Z0Yb;U]1:TUdWCM_V[\Df<:M\N29>4_,03.RZM(#-4FJ>21bM@9BVB79eA9
T1-a[R5d]1aGF@>Ta-?B0WQ-RU4KM)2=LZV#M&=DA1E255+ASYW<SL+,C?#SFaS]
7Me?)H/)X8S)DC+(<1&eW6\c,1[/BX@F]E8LXK-,P/[0:6^?8;.JZ8Q<UE6/Q;OU
_?40NBXeN6c+HL/;P;aSZ-=<1&EAR[<K(TV<E2B\VN=T@eeJ>E^#c=O9^I41-ZT[
WSK;=dcF,d5EGd7P/+2e,F200HH0.I+]K<f\0HVK?;,L6(44b,fW;C(C;B&;Y2D<
YXW1Hfa0(MV@b,gDfUe=f-=1JBM]c5-(<AEXGL[a=P[2YX^4Wb](_666U5]AY)1d
d[3SN6Qc#YVE[2#T#^PX(#?ONc\>6>_)UJGcbJX/G64dD-.gW;af++]4S41^4^S7
2BY(5-9/4L]gD_<:7bEX@=dD)YCI8eE(:1cTF6+<7MbWKUCeYF+Q@TUD>fR.T=_X
R-=)b#?Q=\2(_Z:Y?;e(7)=T;7_G7ADB?-cMW(C(<W)/??.?Z37K@61+g3ESTTOF
O.B8&6C+)Z#?3g098bTbL4.90#g@3#^/L&&:Q4N<7V(e__\WMG]N4fBgNBERgHG[
O<(\A11>7+R90BAB6E9@EW7Ab(gB/JF9N\N(_?7Z3\DN@PGgc/1?_D:4_GZBZV^A
Q5\^Aa,E\aAV^Z7CQJ=B(VF^Yf=R4Od[1P[<dW?BPDY<A\MaSAFd:?\?3_ECR/?C
6R2#R;T3_7C/(0^fX1dLAfZ75_1T&[=+,H;R:BK=e)_:gb?A5JBU]<C#3b&F.<Fg
)E2#E):1+G5]#cT\6]4B4R[HOUaM,GHRZfK&67XQeHC8H78(,8c()\<.OX>/LU=\
bLEYF;DE9)a]_2X6U?9bK>([U95X@)aT[A?N2;a#bWG6A)D0Y&T0_6--XG:[X&AQ
39I0C46_;O3?,::Z(Td]T>?#^V24G7YfVEQ5_@D-=(JMQ=f;+PDa(8M^W>0]-,<f
&aALWTUU#4]M+1E8L0I=.Yb5;3FWd1,E,WVF@J._-SSagSPfFQ.-,38ODGaOI;L]
34FGG\5cI?>0<+@J3WR0Le(5f<\B<Zac^JP&c8/eCOYE=GCCA/?K?KMV#U#@_^@1
G>QT>79I0b6H]a#C?5dOaLad-a3VA^23TR3L_-AfSc_8M,c4d3282Ne\g8[2<[[=
<YFDUD,IH[>R2-LLeeU>MTR;R/-+XZ74S#.)Z5gdD#R^M1:H(\UHeW&E=;.;ULIT
ed_\WCJ5W3@LKB:RW-./VT[eKH_\1U>R@c6PLRWg;P>76DKP)Q2GHPG\eXUR3(OA
H;WAUdIFR\DKN=NQ\\[@PE1c4RDPG-PW=U.TET,]VKCASf&R2BSG\0V=OdBKM#W_
7(-dO_EKCGVSWfa+F].DeW33b6XSY?D8:dbK245#aF7H[4.F3:g6I)^)FJ[42]\:
]XFY44<#P+;^WHDF1\FP/K0WEWKgVNgcV(QM5TX#eEQ)LEbK+@RBbS6@I+[CI]K>
]g>V2>=[8@<g8)-#S?>^1;9K<4:=5&5L--d#:)A<G/6=+Vc7Y):8K:;\EEWEcRg]
SN5bG,gA\1Mb:[cO^+W7+=YDHDVCPS/@D2.[&=aDR5&X_(aR2gQ8_bTQU.GL@Sf4
W9M?N]M\A+L^FITOXH.9KF[GaH&7GAI.0/UVS@I1KT6)31QCPRfBH@Y:J?3K/30B
<X\PY<U1g(UN#cE)ef-5+Q9:dDTL5M4b)<LOZB?B:X+>(dW)U718Cb7/=W#,J9_G
[82N4K[7a^4L6959(-#O#>.II09>B=>KbOF-S6a+bFW@#L+1_/8&M_9e3BYYS4QT
]bZ4Q<<EDNE^\M\Pbb4Fc7ET.b>Acg5.NGM83S#6+SW7+KG1EO\.&N7.MZb,^E,e
GFM,8-UH7&IN6UeS>-YZV+_OZ#/67D^0..N+Q3\gHEgA:AXeQY/.d<0_+#ROE_R2
WTX:d#U#[0JQ&LKF,-f7g()aODK7;SfIT4M9IND[>K\YQU;@Y._0WbS/8A?8UV&(
&b@]-cL#df#NLH#eY#9M8<UZY0YDdg-#be]#@,C:-a5[IeQbUP71N789;_D=:]ZO
70&ISW,]-S]7&4SSDWPdE@V,_0Q6[@_af+]5W9HK1fc7YS<c.bWFTWH&d#MZT2G)
NZPKXF1e=&=A+K32MJ[c,+dU(G;]8;E)b2&Y)EKNT3A_Z&VRa:3QM8F_PAa8E5-@
:3gFX&f=1#+MLbNJV\6AgP7I?)F[FKOECO#J9V:UWXPTCP+6_L>I]8JYGAN2(JCb
O^WJ+HfU^WYd@3B-Aa?4747_f^4VLE2O6YUgS^)(R#=a\PX[/A]#Y(\>e<TOd6<&
B+J&CL)63aPdc3g@)@N@@=L-S4;fVB12.2]&RFMF2AGI>@WW>[<LUW.3UX&,0UaX
c@K>E<RC\&N+OI>E7P2\)HbNNL1FJBVU67/S]2<3Dd._X^^\RZO6VX.aPa5T\[#]
_fFI,XUWd5-YT[VG37Y?g;U<)X1>9g+4.J[4E#T&?YN3Re(.<>,1cS)J#,CB<^La
aS72W(83)0MJ51IY.dYbC;#^M.eC@&C@4.5K^)+Q#4],P=9L:_Q:,WFgCaR0H_+N
6<D0bS38P\XILF?FS4P&Cc+W0?LT5SVH)FL2XVW[6Ta.3ZWGP7=H:]N;M:eCW/eO
+E[BPO5Rf[gSZ12:fbAQGA/^W:]C@QBF)Q)[5BJ#>7;5cB&6GDB9:G^>IKTH2E[(
eU5fa9>\@VX1V1M[#N;D23M:fLFF;]=6-5)_KK.HQ\[;EWaYR\&f49P_7R>?O&b?
5D1V_8;eTQ8K>6VW[HSB/LA6RAV<)BG/[5G#8=J#cbLR<TS;W?<c;_,N]VbLY/4a
fQ4J4(1<Q[D2^\7-A(^7,/N#]C3_J@+,^,9))FPCQS(Y7UEN7(#&05de#G.NaegS
R&\=.F=VI^/1=S\(APKEcc<fcD84QDDgX;>2ZG_P.+VS_]JN_SF#f@:dU,4X1N<>
>_;ZHY->-)L=^4H\C#BM;XLX0;,.11X]#S;W^=:P,LJ[VS26L1JZHB5_-76;f>96
1PAf:X=7L6b1@+Y>-I#\N@M21A/+2\H2O7VWLUG05=:AR3YDdY>=DPJW_]_A67V/
PSRY&-&,@0HSOQ+I^5Y_67Xa;LZ0J:MRbI&[0#QN8Lf#30M?HfgFa[:&]TYG\2K4
>fK?TP],U3V:N+[V:#_E@2]e^b3[F.ff&R9B@90>2W.S)?BYFM5AQN#4F(Z8?+J2
(5a&Mbb5KV6IeI?\DFSNf.JX@,(I&N&aOH]G/B-_Z3Z7g_9=&C<E&C+YMW?E7e_:
<K=WHEG6#WNSS7Rdca]M_X,V)9(2782R-<.aFX?Ig2KI_8LZJAA(E&>Pf&QXHbJX
BFAAY^V0-W9D&=D\\ABDcP3E-f:N&&cdeH]8>?HKSW?fD-LFfLS]+b7g0,&f.3b<
F-aC7[KVDJ2D52-H-GYO;>]+<)KFCAL[f=>C-X(XS?.C5.Kd,.A12WQQ7+#bTa&A
,#@MgC.G[D]=36YGK4=NJ1,1VY.DX@0Va=IOCLf7<PRJ=dSL>3/GHW]Hg;C.cCba
/<DK.]bZYQGf^<2f(YP2@5XRb;@\R7B#ePUP7ZZ:5@\b:\VELXO(CB.>2&8>K>^Z
V_FO2O<\D<2#fQRSYFb/>eW-BfRe?WI<Qf=X\gOca]#GMaX94#(6U/N6]<3UMZ]S
E]..8b\GR?1\B3Cg=[/9>DV88=8aVMS-O#HKa8=gLI_R8HZ09Ec^DQdD[(K;5@K+
8)KcT=JYLBbNbVf(T+Q?T&MXKNLIIM5@cEXFbd).eQV3N-6R<57<-X9#=-2;?[3I
gcA@Yf.9bbOT7#1B1d&(;Q:&SE:R+;@]/+3JHb7)=4W3Ig<Jf51/+fQUHg:O83ba
geFOT>5L?b@6g=[c_?9WRS)<PZ-[HO#=_5D/]93?R2g:aVMbBKKK582:VNZ<]T@>
.g>^d75_N?8&-=E=Fa_GYEHMSRZ;J-Y,U79WXNYV)Z/+2^TOEV-caI,,(R/fPDMK
02aUg]W\5LOJ66@e<OSf/[,(_;WfS?1A+T2CF@d34K_f>J(6D=BH\Z]_T]2Td-P9
g@AY(8N.JZ04+<828VQ2UXSCARC.F#.eDM\,&/2,^PZU61/7]S,=b,2YJNfCK75e
c]R[^D-)EF?T4HLI].RL;HQ-=)fc(S39<MTH]-b<VE/333MGbID&f4TVaM@LAKcS
SfM8Y@CSHXKQ[b>GaUBVAY:ZV94\SU-;Q&_Z4Y?3JKUZN216M;f5YWB7D,-HgUK&
UGVY00<=BM)&4V9E2:?^9G:=_eK[MS2>b-\L_TK&QJ;Kb_;a,eG4VF=AXJ5\(07D
#0#SAJJC@H3;JbOW[)X,/T(-X^H_S)CHX0VbZ=].&e7]M8D[855K_UB29f-7.Q)A
:.d-2#JEX-ZQRHOR6#M4gT/[\KB@?cJ^4_O&<5VXKS;5GUA,S:9Z0D)RVNOVTbF/
ZUZd,]J+g=cDc^#b_MaaaeGV=]&D.)>a+.]#L7V)#)^?Ba]R_Gc^\SV0gT)&Q7V[
#D<X)W==D(=eSM:Xb5>UP\WW.I;5[ZI:;Ugd^FD;O3:1Y:@g&0bY0J?347d^Q1[B
>[@W+77WH/OJ&)RF(5dMQW.LB.&G#6FB^2IECa<.]c.?].S.cHR7b7f-BS0NJZIR
Ge/gI.,J[gP(Iba87W]BY>]#M\Ne,00?@EV=K=,g(ca=cMAdC(aF3XF3GY:C(AJa
6YL>0G.0U?U=54@@Y)4_[0\>,S?N<B,P4V5B;+CZb5(:J9U;W8KcRNWCH>0Ic43?
WZOc/:+37R#R5]_MW4;g=(Sb+155KUD^SIc&XJ(AXa?WUFJUEM@B3LVf0,eJ(Q>5
KVFL2E#UR^-JA6E_IXa][JJ9S]XP^&G.E@3]bA3YLS^N>Mg@M;/=MKR;K\b^6LgT
Q^@N\I9c6bcJ-0Mb;/7RaZWd/GN#beTCGNS7e+#AWW@\/X<XOcC_Z>)MS]SG;MWJ
?2</UVZ8S6-.CAEgbZKag\B8efYf).JR1IP;\I(35(\0b17\;=;JX7Y>C#HHVW.[
X4&Z4G[OYY/HU@>RU0ES48=._R+@#1JeXFgHZE/_e@&Md[c[@1>TfWIIB\XYVH(2
Da47gL9g@(dPY&CL@g,c/<Z[]N^[8c:4SOGSG65.N/27M-AXeL-UXP4_X(;^_Jf.
=_Jb6KDWMP?6C7++eQZE:3W\E-K<&UC/dEX(+ORT5//J.LfEdg^?ON4H&dUVP9K.
G87HgTH[O#AT@a0f.Qd_Z&Z[W-f:g,>0HIH(3EGcT0L<30gN:]A(/\ALEf409Y3g
;P]K/-M^>?RZN]A44_KCV&(7)#.L=0P>E,\.?f:(<\E:E.BH:&E1\/].7>.FGSL-
Oc2O7gdN^B2d],D_]aCK)VI8;MY+\=E.QTAd\M)\EK4G=3Z,8+7=XRBF3b?GU9TG
F\X)@K?Y2S+bTABT,-L]CT,S\8C29c1_0FJ?N22\)a;d,^]a_a-c=XB0_QE+RLOT
A5B^RUA6&?-D-d<9(=OafEC\HdG]884g(B<UJXd(=5JK471.bCK-LK&/-ETc,?-T
AM7AdUgQ-dEd/,QUU6D&8>#9JM2KP(3X(^A9bc.GYGPbL.[7FX6>4E0P[1IEcE[H
CHdS[5a.B?B2D?6GbOfY:bLYV6G)9V1TXf._8SE7/FPf8beceLWS/S1F@-](Qg&,
Qb:,Y)_^SgSD0O\.[G)[gHXXL^Sc?W,>W_>EENCaS(H0DKG;ASA,MgN,(bS2E145
L&X&MRJ#HRJI]@-R+a2&BT^OA:5+c(EEP;?9K>?XI?<]]P6T)B-:/1aQ:[N@XDaA
#\V29DMZ7f+Ua^^LNeAXD6[C@=,LK7M^A<Q02/7R<1+a\--RS94_)]QL&KHJ4OH=
PDU73@BeC7SVT8A&:D1d?IB9H+^\J4/W48C@GR6=b\?g;G0E;HY?BRPRJ_<9E&Td
AX3PU>#.-U8HB;Y\#4H-=ZN4W,L&\S9-QVGG;55bF1ICEQe;QXF[\K0W<CZWD\@3
JA>[Oa-a3fM.A9OBI]FG3^ZeWSg_BY(?>Z:LTW4H<R;H=[4?;@2G=O]KKcTR@d9I
[OIEHe[T?;VPJ@7>DK27WZ;GK^?)D^JGDc9?\DcQ5&P5Z_.C8D+>61[AgZI&,ea0
Ae;a[B;1K-O3GTa-,=O<?]fN7M8ZAd]9fcOMSNfSJ<DK2H9+JE\1XN,&Y-&U[)fL
K/#3\Q:N>B)=H1:1UQ554dRAZLbRaEJdN[FI1A:AcVN;.;\SS,>(M5@(#,ZX/1F@
O2]<=>Q;\bX.)]TTYc7VHDaE5,C>B4S9<A&XV5c6?QZ+C]Ge5c6NO&3TAZ]<&LB]
c>DH7ZA6Ie81F-,BG(d^(M2;[C\83aYe4QZH8)P+BWFLa[bZLHA\Q/]2G<W..::V
\WcXV7/GTKH&2-7@eQ/82d>bGNP=fDHaEd6MX=531&UZ/8d@cc>Mc-/5S;[<Fg[,
D<5\=D;EbaD<.f&;M8[AJ#+BGd=/P^aQUAHTZ7Wd&fLG5@O+64][a;BcI7ULREDP
>+OL^B5+aF<C5?:CaG&8XW-=\NMV-JNK/GN9-BOS5B^[N>V/]#4K0g&+DPA5T9Ia
3X[J(XA=.+9aQ9(XG7RagMa:9I5MgL=4XTd&+;<&JX8-6FUMc5GSA_M_7_<D/OW9
(W[c<Y0<cI2??f4.bgS06MV<BP(QB>5<;&O\T924[C0QS)B)eQ6Y1:Q==+])QJa7
CBB^MX\8_SfEV)M0<K)CRedE]\@UcCb5B5Q)dKXI&&QDbFJcVRQ4QE^]7G;/Yd^e
@SScLS9GdQX1(&_O@1?5UT5ObF85ZOS?@AA&fSQc0FYI/T_L3(?W[a<.#J#LEaFV
bE\.KG?76-\MJPE08C1H3/>T1BREXI?K4#3XgGC?D4K1GIFR\TXc)@#(aS6Ceg3a
A7c2^;dDN>)D+EI?6MIWC&:dK3PcI_2Ad>[\2)016-gKJ5^<SC84g=ZD\8VM2c1B
FT797OD_T69L?SALF65:2a[^Ua7BYOX]cOFJ7@,6IZcJ/E3E^@O/>WGE>]FM5\Q;
X0)1MW5R?.@ff(WN0H2L@U4>6aO,J8<:W5HbJAJW]EO2A0:K7]gTQBT87Y1e_C)]
:B^GX-C.6(&-Q?._6[VNWe8YR79)8(L4G#dOE\5<&;3cV.a2[=]b)#M-EeU8RdT3
XdM&f?V:b[2\HR9DQYfL;C2CKJ?0Vfg4(@WFY75X[caCd>2=MF(4[33?YSG^5R8K
)B;fHDgdG\10\F\[^e\/9E?VCa?f\JE#6H78+-8[K@@-g.KN)/LIe.7^M67^E5Z^
7<Tc_NJ,1S5@/bJV0JQ^^[CKRQb4](;]MAdIAZB65K-OMe+T+EgV<T+f7,ZZ7WQ<
<2ZP?<7baXVCKaNI)bN\\UA/LXVA4?]JH:-VG6PQY36ZeP1I3LT+(Ob:.Y]H8HbL
ZF#];H:.>-U)CUcKW;__.NWbN3QP),18<b&0\Mag7_;Yffe<#RIM:B\&35XWX36A
F2@5eSG@5,fE90D82IfN,d+\,>^EQHDBM)T#IJ&FLMee(F1]S+NY<f/<P#7[TCAH
0S:95fNS7E<1O@GH?7c^OQfEeH0;\.Sb]8=B>c96K[9T3,^;,&29:AEa[c#,(ETQ
]UUXMIE8ZASf0_YI\2PM#M(/H?>g=?#Q]7BZ<,>DF.cd<.[W.B.@;S6,)&X#(#8L
Ma\Z&SY\;LB)+-cJ3O8APbK(2<4Ce]P]?V]3be3S[D7]BY3G>>LLf,&V;I0GI+[=
5SNARO^#J7c3H?7d#GcNNQGdZdN\,R>NA,,4X&/FL:J0bf7AA@M7^MWg=GIZ)KV/
LR3N6=(7MHGe.,8WYF[;<QY/P>J/=09Jg,]AG27V<H905OI_+CX-&B<8JMa1(QXD
N#C-dIaXa2;OD6O:[_Z^\JS[aK9PW4?:V;Z[4[ab^V9XL8:E4=?)LPG7N(^a_7aS
6L4G?G6U(0gCRR.C3UQONc)1&9RW0D_5d]2W0UULD&cT4?<7V0(I#g1a[ZZ0JX(Q
CZZ3KdQ>5a1,[ECe>DQ_@VDS[[ZT-V6BgB3:Y?c=+9F,:be9I\PU#Q2&+77U0K1]
^agG-^NOD^\J7)E/O+0F6&1=AKD7@2Pe57&e&aGcW[L+/83BWII_Q^b8JCU2gPJ0
>X/d85KU67(^(S7@YE6dDZK0cRWMC5fQSe]#b.@F(WWQ+-,g/BF+\e[93(M_2GLA
9-.3@=#<DFJ6_N<YX)?++DT@-4.([3YYTC[d3MLPOJ^-J)^-6:9,L.g9cX/=-BO7
NN[I@8Y415WcRL0a,&7XO--0CPAZ8\PT^Z(DUf8V)U+?+/IH_UbVTJ4.-3,#C^.9
^Pf:6-1;A6[_2M&CQ(#>Q0PHSg4FfFS=BC;FWL=LIb?A029JX0].EdcJd/<geU(M
DNKbGeK+.ARce^<U=>4H]C<[(&R769-ROEB_J(4P(6)EFE=cg@6U<+Y=+/UBAW95
WEeK5HIe+KQ(2a^@]+16J(^1,BN5G(2-MfUfW7f(;P(IE-B:49]^d_gI]\&<[-8D
MbQ9:KDA)S>GL/T^df5,_]C0DK:G9dDC8]Y0K6cZ>Bd7MSNF9ST_2>RXZ&(J5WcD
.#^;NF-e6T<MKaeSRO?5IBfXd>/cb,,6HP43DD:7LO,S)=+&)1++b:POQbLd=c[9
<&@>:?BOJ;8FI4@>OP_#]2E)58EV\?]4:5._D0WV(B/X=X&c(E/.N/<):H^VYQ\a
P@acB:@ZR-6=8dgHe^ae\fR6R3]LJ816W8\_gRG?/0F]\KG8Yb,[^b_4a\[UKPR&
.<bXeJ]W)LFH,LF>X]N_8(Fe+0^e:BC6(KY@+Sb>LXR7M.LG76D<7S([;YbH2>B(
NgF27f8&-#dQ>93b=fLGQ26VRWFE)7M-f,MR7<9,;@aUKC,>0-S+H11@<SNW>;F8
Da7:6FFK3OK@)60a95?Q<RU^aH3:5QXMWI,#F@aVafO;bCDBbS4^]&,d>FSb,b;Z
Z&]G.>BRF3RbR-ZQffWYdZN]QEZAE4;P0JQZ?,U8M3OUO03@C=0I@D7d0/GAbW@F
FW\S5daTIFF+#Sg>\[L4-+c73X,?I6@AQMeNd/:?3A<S;-+52Q9UJX>=)dI8MVT0
2&W24Y(45fgD6C5dd(N/-0(.f#U#E@Sea[RSbSWT^^7SR@3X:\;7Q@1<#JU9Z[^L
RN1)VZ]Y/dZUAGbU.@]H3bHc[FeHDR7COT[.5.Gf&QPW1DfS]7NW6#/T+fPX9Ad[
<NL2)>#Ze=AdYO;Y<HJ1b,aX5QPLNT]7.K37XM:SYaAdV_P+O,/<VMOfWeA\-B6,
NKafZEH5W8<S:Lg@X33?JFUc);bfA2^YOCAW:;ZS:H:g27SZ,=5Z[-b7bY#I)2E+
=;N5IH]7)d-(,KbNB>4?1+UX,LH;B\d<X,_J[c-=@J[dS:DK.IOX@LaC6e+eM[?:
YWGRDaT^0)EcK&(e1IT8T2025-&RN<8DW@4Df:D)R1gJETK/H1SS]6R\+D^07.Z)
6IRTg,.bX=LGL(GF96I<;JbAT1RW(DK>/V1eHVR0N)##K7.DK388,=&-_QV#IM^P
8B>1RFQF=Y+BD;(:_0OBb:S6JZ.B9)+H&CH682.aff/6[.239SEgg6,X@:TCB+S2
)fEcH.Q3ISCA:=-ARZ1U#gL/^2E(bN0G[+GGG&9+_A<:@[c/D(L>H?c+_I/(BA\Z
91K0MR=R?NC[A#gg:EbTG<4+SWW:PcD<EZ#?aQNEP62>E,\2LNDER@4S^G:Te>TF
M]4D\J/C4fNB:8-@?H#HQ=>MYD=g])W3[5F>eE(G(2:Z.BV/IcS6Wd?I/8dB>:Xg
Q=W[5+P9B5^7XKAW>@,;d&\<3[&^K^d9bA#1D<C?eT[NaW\YQBc^J5^T8=R<VOI+
Ffa&Y?,5f,XA023R,Yd8\aA8F(DDgeT9K>DG.;OO:5<X1aZ554#0RC_RfE&4Yd1=
XJIBY+@N;QVXB>.IJMZOT>d9SJ-2G52NG?F<2ZEXRe2bG(E]XL?a+c6@O,WL3=OO
V>S.J[.3^K<[:&8XfVZ/3BJC@TT&bZab,446#IHU9N_Y14=g\a7[dEP[LV[=-&&@
ZMBYG^9V-77/@fHgVOYYe7F?NI6W6+(+^U6QE#aKb#;eZV[#-\9@aL:gSb26\g[6
5U3D^JD6_][9RQFM6I>H71@EV\\VCgD[>4eZP3g<;K3I7-bd)@gcPIEegH5NC+D9
9BOfTILEP<1:UQeB(0IN,\Oc2LL6+SeCe>@]=)Q)7:N5#+KUACU8,AaL,EHHUN4C
6#eQ6TEf#0DBe;.#b>9L2Z<7?5gDX#&JHSJ0L\\42<E+3N;Z,M[FR:Y@)XOMMcWb
BXCPMc-<>IS.^Z5F5<WSZXGMO>]O(BLOM;KfTgCH]<=fSe?6CG5a_6dVgB:NC53O
UUU;0eYbZBH]^&0R;NA((WI9XMBe(EcBCeN4C[^#@?fS@/<GAV_6(QN.eD6+=&(?
g\_Z[\9F3=1EC4(gO_WFcH1ZT]7?,=@C(@>T3<&]6208Y#S15.g&9<;>gaV]e7E)
H?91bQU,@:7NI\HPeQa.STb@3)578J;H6&ATP?HH,N<QFE77,393\]LJ>?]6USU&
2&BNQ4[[4#NQEL:5eGV)]<\VJXBR,?E-?<S4c>RM1;:ETTO\65K<.eeV=/3Lc=D5
\V,9Q](TE5T&O7;;T8^)7YdDKQ<BD#\2:@2eL39#;.VD^:\4>6Q<_eA[Ia\TM6(9
-Yb.-MIKHcXLO#_=A5R#)WV3;JXKeF&4a7O#INB[5_(c;D#MU#U>6H^MB;4BgP?g
R=Pc_.Y_AG7DXH5&e/dBPZHR+KB-#IK51db+F[^3Q8B:AC\Q<YW[2QHD30,F7bG4
A;6/8DWcg3,A_>Y<[c_GgZIW5:JQ3Bd>FW>]NNe<A95P/[@JEK_VU2K2+IHY&9A_
,EbC<S41XB;AO@7/8MX1#db6^.XM0]fN?/5(VWaADT5@=4)-IHVa#D3/M@&bT@JF
8/c=SHHSPgI\#K[]KR2_HV)@X=#)=HI\8R;#_5PI)&C)VVLcf73W@[&A6+fL^VL\
IebFE:/=\FX5bD/16<>IPZ3g=L((UXQ/M2,&6;HcT=GPg02G4V3^^<a=7?eD;>1d
#EYbS)MV8,3C8G[1e]AHD-K)&GETdg\gc=1K@UB>KIXIcM4@_Q9/7;ffH:@1\7)1
dH?LE>WId)_NY]aOS=LTEWf_(A/baN,--YT2X(V#RIL2<I#NNcS\e,WdJBPcG#>a
G_]gABTP)cE#ZbUb,5J=^G9^L37#O.&@7Tb-S85W_8?dLCGT9DG-])ELJ8D^NRJI
cf-)J5PUX5164-:=TU(8bOA46N<dF3I8W/)NIS3,W/@=:)G;#??:geUcOLIaP:1[
(<b]/JEY.UHHR^-[g/6K5ePV1K6.Yc=_6+(P3-X)Y^DQ=DN)],FCCTPe[RCQ>IWP
V,4)L6T=\,FU?RLbK]J9)M;,9d<HUZ?3F)U^V1.YOC)e9dJcRQ4&()0f,=3J_B[4
A@C(Q5CFBLMX03NZ]_XD<?[#1f1EJ2dgB;Kd7>@c^GB4,>OH5dKTO3\JVeZ;?),X
6E5OB[Ya.N[TT?]D<8UL^3.PeZ1TX&I77PD0g_XISK1SNGBbCc]/TY(V?e\J,MQ?
^L^282;\(6Sf84(>M3f(N-;d4_He8<YXRMC(dNMS^WC;YP4+N<S:UT+-.]:5^]Ka
Y-CB3<:.-_c&F5d9S+</.A\3B\Q;QAV?.a9VDZP1B[8OHP5bZ-2@B2A]D&_cED:V
UZH[U=>/,EcAdJZV<>UGc^f_MPZ[5SR+c7EefdQW:>U0>Z@-Z)6G^HROOD;)[(D-
T?2dbUU)>,#eJg2G/GCJT2+6[:V[2#I8BgO2KF4S.6NJZGe/Q[;/YJdfDF=Z[cCA
X93@a@=W4:>FO,D]6@/I7J^@N.E@:f6WBW,]TQ>)7g,>Q<CJLbYU3A^6eZJFQcJ_
H#(/@HN?P?f]66Q:NfAP/;+b=(/8e]YWNRLAYEeS+cf30_6f+IEdBET4IdST>S41
T[_::<94G3P&P@3AV=<O8PO4bKW.E],4U3VCWN),OA@ed0TG8#RNZT33a<HRC?DB
/23F+?M2E?RJ\Db?]+&SSJ06AIT/cGC;8&C9-LGJ_DAcPTTKSQc/3)KN[Y/3UM[a
SVf19]RbB]+\a8e28Q-#F]X[](\\YP(B_\bHEe?+SW6LZJ.8S(ZCE3P-D:^QTTQ5
^(D,8<2;a3#+F5FT-dB#08bO87@NKLF/D+B=)_+gOG311.@f#7^5Ab@8caW)I+_W
L[:L#W#0&1R-AKRBVGX](:;C7ZU31+/B664<(=2-WV=I[L<^=[;B[48ZO/_(2XX0
<W7JIK]LN@3NUMTC1<+GU]664aWZ]ZJbVeCc5&N>\X@UYAV[cUYc:0)M5;SB3@Y(
))]ROgE&PdUF6Ka_N=1NMe6>OXd-M=IC=@b4-:RbI=S](F&?;J)RJ])ML$
`endprotected
endmodule



